//version : v0p2
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AD1HDV1 ( CO, S, A, B, CI, VDD, VSS); 
input A, B, CI;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B, CI );
  and I1(a_and_b, A, B );
  and I2(a_and_ci, A, CI );
  and I3(b_and_ci, B, CI );
  or  I4(CO_temp, a_and_b, a_and_ci, b_and_ci );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AD1HDV1C ( CO, S, A, B, CI, VDD, VSS); 
input A, B, CI;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B, CI );
  and I1(a_and_b, A, B );
  and I2(a_and_ci, A, CI );
  and I3(b_and_ci, B, CI );
  or  I4(CO_temp, a_and_b, a_and_ci, b_and_ci );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AD1HDV2 ( CO, S, A, B, CI, VDD, VSS); 
input A, B, CI;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B, CI );
  and I1(a_and_b, A, B );
  and I2(a_and_ci, A, CI );
  and I3(b_and_ci, B, CI );
  or  I4(CO_temp, a_and_b, a_and_ci, b_and_ci );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AD1HDV2C ( CO, S, A, B, CI, VDD, VSS); 
input A, B, CI;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B, CI );
  and I1(a_and_b, A, B );
  and I2(a_and_ci, A, CI );
  and I3(b_and_ci, B, CI );
  or  I4(CO_temp, a_and_b, a_and_ci, b_and_ci );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AD1HDV4 ( CO, S, A, B, CI, VDD, VSS); 
input A, B, CI;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B, CI );
  and I1(a_and_b, A, B );
  and I2(a_and_ci, A, CI );
  and I3(b_and_ci, B, CI );
  or  I4(CO_temp, a_and_b, a_and_ci, b_and_ci );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AD1HDV4C ( CO, S, A, B, CI, VDD, VSS); 
input A, B, CI;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B, CI );
  and I1(a_and_b, A, B );
  and I2(a_and_ci, A, CI );
  and I3(b_and_ci, B, CI );
  or  I4(CO_temp, a_and_b, a_and_ci, b_and_ci );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AD1HDVL ( CO, S, A, B, CI, VDD, VSS); 
input A, B, CI;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B, CI );
  and I1(a_and_b, A, B );
  and I2(a_and_ci, A, CI );
  and I3(b_and_ci, B, CI );
  or  I4(CO_temp, a_and_b, a_and_ci, b_and_ci );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AD1HDVLC ( CO, S, A, B, CI, VDD, VSS); 
input A, B, CI;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B, CI );
  and I1(a_and_b, A, B );
  and I2(a_and_ci, A, CI );
  and I3(b_and_ci, B, CI );
  or  I4(CO_temp, a_and_b, a_and_ci, b_and_ci );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> CO 
	 (CI => CO) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b0 && CI===1'b0) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(B===1'b1 && CI===1'b1) 
	// arc A --> S 
	 (A => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && CI===1'b0) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b1 && CI===1'b1) 
	// arc B --> S 
	 (B => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b0) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b1) 
	// arc CI --> S 
	 (CI => S) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module ADH1HDV1 ( CO, S, A, B, VDD, VSS); 
input A, B;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B );
  and I1(CO_temp, A, B );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	// arc posedge A --> (S:A) 
	 (posedge A => (S:A)) = (1.0,1.0); 
 
	// arc negedge A --> (S:A) 
	 (negedge A => (S:A)) = (1.0,1.0); 
 
	// arc posedge B --> (S:B) 
	 (posedge B => (S:B)) = (1.0,1.0); 
 
	// arc negedge B --> (S:B) 
	 (negedge B => (S:B)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module ADH1HDV1C ( CO, S, A, B, VDD, VSS); 
input A, B;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B );
  and I1(CO_temp, A, B );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	// arc posedge A --> (S:A) 
	 (posedge A => (S:A)) = (1.0,1.0); 
 
	// arc negedge A --> (S:A) 
	 (negedge A => (S:A)) = (1.0,1.0); 
 
	// arc posedge B --> (S:B) 
	 (posedge B => (S:B)) = (1.0,1.0); 
 
	// arc negedge B --> (S:B) 
	 (negedge B => (S:B)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module ADH1HDV2 ( CO, S, A, B, VDD, VSS); 
input A, B;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B );
  and I1(CO_temp, A, B );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	// arc posedge A --> (S:A) 
	 (posedge A => (S:A)) = (1.0,1.0); 
 
	// arc negedge A --> (S:A) 
	 (negedge A => (S:A)) = (1.0,1.0); 
 
	// arc posedge B --> (S:B) 
	 (posedge B => (S:B)) = (1.0,1.0); 
 
	// arc negedge B --> (S:B) 
	 (negedge B => (S:B)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module ADH1HDV2C ( CO, S, A, B, VDD, VSS); 
input A, B;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B );
  and I1(CO_temp, A, B );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	// arc posedge A --> (S:A) 
	 (posedge A => (S:A)) = (1.0,1.0); 
 
	// arc negedge A --> (S:A) 
	 (negedge A => (S:A)) = (1.0,1.0); 
 
	// arc posedge B --> (S:B) 
	 (posedge B => (S:B)) = (1.0,1.0); 
 
	// arc negedge B --> (S:B) 
	 (negedge B => (S:B)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module ADH1HDV4 ( CO, S, A, B, VDD, VSS); 
input A, B;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B );
  and I1(CO_temp, A, B );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	// arc posedge A --> (S:A) 
	 (posedge A => (S:A)) = (1.0,1.0); 
 
	// arc negedge A --> (S:A) 
	 (negedge A => (S:A)) = (1.0,1.0); 
 
	// arc posedge B --> (S:B) 
	 (posedge B => (S:B)) = (1.0,1.0); 
 
	// arc negedge B --> (S:B) 
	 (negedge B => (S:B)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module ADH1HDV4C ( CO, S, A, B, VDD, VSS); 
input A, B;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B );
  and I1(CO_temp, A, B );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	// arc posedge A --> (S:A) 
	 (posedge A => (S:A)) = (1.0,1.0); 
 
	// arc negedge A --> (S:A) 
	 (negedge A => (S:A)) = (1.0,1.0); 
 
	// arc posedge B --> (S:B) 
	 (posedge B => (S:B)) = (1.0,1.0); 
 
	// arc negedge B --> (S:B) 
	 (negedge B => (S:B)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module ADH1HDVL ( CO, S, A, B, VDD, VSS); 
input A, B;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B );
  and I1(CO_temp, A, B );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	// arc posedge A --> (S:A) 
	 (posedge A => (S:A)) = (1.0,1.0); 
 
	// arc negedge A --> (S:A) 
	 (negedge A => (S:A)) = (1.0,1.0); 
 
	// arc posedge B --> (S:B) 
	 (posedge B => (S:B)) = (1.0,1.0); 
 
	// arc negedge B --> (S:B) 
	 (negedge B => (S:B)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module ADH1HDVLC ( CO, S, A, B, VDD, VSS); 
input A, B;
inout VDD, VSS;
output CO, S;
wire CO_temp;
wire S_temp;

  xor I0(S_temp, A, B );
  and I1(CO_temp, A, B );
  assign CO = ((VDD === 1'b1) && (VSS === 1'b0)) ? CO_temp : 1'bx;
  assign S = ((VDD === 1'b1) && (VSS === 1'b0)) ? S_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A --> CO 
	 (A => CO) = (1.0,1.0); 
 
	// arc B --> CO 
	 (B => CO) = (1.0,1.0); 
 
	// arc posedge A --> (S:A) 
	 (posedge A => (S:A)) = (1.0,1.0); 
 
	// arc negedge A --> (S:A) 
	 (negedge A => (S:A)) = (1.0,1.0); 
 
	// arc posedge B --> (S:B) 
	 (posedge B => (S:B)) = (1.0,1.0); 
 
	// arc negedge B --> (S:B) 
	 (negedge B => (S:B)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV0 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV1 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV12 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV12RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV16 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV16RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV1RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV2 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV2RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV4 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV4RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV6 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV6RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV8 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDV8RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND2HDVL ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV0 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV1 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV12 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV12RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV1RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV2 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV2RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV4 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV4RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV6 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV6RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV8 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDV8RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND3HDVL ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND4HDV0 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3, A4 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND4HDV1 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3, A4 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND4HDV2 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3, A4 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND4HDV4 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3, A4 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND4HDV8 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3, A4 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AND4HDVL ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

  and (Z_temp, A1, A2, A3, A4 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO211HDV0 ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    or I1(Z_temp, B, C, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO211HDV1 ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    or I1(Z_temp, B, C, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO211HDV2 ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    or I1(Z_temp, B, C, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO211HDV4 ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    or I1(Z_temp, B, C, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO211HDVL ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    or I1(Z_temp, B, C, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO21HDV0 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    buf I1(OUT1, B );
    or I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO21HDV1 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    buf I1(OUT1, B );
    or I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO21HDV2 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    buf I1(OUT1, B );
    or I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO21HDV4 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    buf I1(OUT1, B );
    or I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO21HDV8 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    buf I1(OUT1, B );
    or I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO21HDVL ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    and I0(OUT0, A1, A2 );
    buf I1(OUT1, B );
    or I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO221HDV0 ( Z, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, C, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO221HDV1 ( Z, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, C, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO221HDV2 ( Z, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, C, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO221HDV4 ( Z, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, C, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO222HDV0 ( Z, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   and I2(OUT2, C1, C2 );
   or  I3(Z_temp, OUT0, OUT1, OUT2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO222HDV1 ( Z, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   and I2(OUT2, C1, C2 );
   or  I3(Z_temp, OUT0, OUT1, OUT2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO222HDV2 ( Z, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   and I2(OUT2, C1, C2 );
   or  I3(Z_temp, OUT0, OUT1, OUT2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO222HDV4 ( Z, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   and I2(OUT2, C1, C2 );
   or  I3(Z_temp, OUT0, OUT1, OUT2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22HDV0 ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22HDV1 ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22HDV2 ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22HDV4 ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO22HDVL ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2 );
   and I1(OUT1, B1, B2 );
   or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO31HDV0 ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2, A3 );
   or  I1(Z_temp, B, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO31HDV1 ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2, A3 );
   or  I1(Z_temp, B, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO31HDV2 ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2, A3 );
   or  I1(Z_temp, B, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO31HDV4 ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2, A3 );
   or  I1(Z_temp, B, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO31HDVL ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

   and I0(OUT0, A1, A2, A3 );
   or  I1(Z_temp, B, OUT0 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO32HDV0 ( Z, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  and I0(OUT0, A1, A2, A3 );
  and I1(OUT1, B1, B2 );
  or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO32HDV1 ( Z, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  and I0(OUT0, A1, A2, A3 );
  and I1(OUT1, B1, B2 );
  or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO32HDV2 ( Z, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  and I0(OUT0, A1, A2, A3 );
  and I1(OUT1, B1, B2 );
  or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO32HDV4 ( Z, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  and I0(OUT0, A1, A2, A3 );
  and I1(OUT1, B1, B2 );
  or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO33HDV0 ( Z, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and I0(OUT0, A1, A2, A3 );
  and I1(OUT1, B1, B2, B3 );
  or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO33HDV1 ( Z, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and I0(OUT0, A1, A2, A3 );
  and I1(OUT1, B1, B2, B3 );
  or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO33HDV2 ( Z, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and I0(OUT0, A1, A2, A3 );
  and I1(OUT1, B1, B2, B3 );
  or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AO33HDV4 ( Z, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output Z;
wire Z_temp;

  and I0(OUT0, A1, A2, A3 );
  and I1(OUT1, B1, B2, B3 );
  or  I2(Z_temp, OUT0, OUT1 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOAI211HDV0 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(B_inv, B );
	and SMC_I2(ZN_row1, A1_inv, B_inv );
	not SMC_I3(A2_inv, A2 );
	and SMC_I4(ZN_row2, A2_inv, B_inv );
	not SMC_I5(C_inv, C );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2, C_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOAI211HDV1 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(B_inv, B );
	and SMC_I2(ZN_row1, A1_inv, B_inv );
	not SMC_I3(A2_inv, A2 );
	and SMC_I4(ZN_row2, A2_inv, B_inv );
	not SMC_I5(C_inv, C );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2, C_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOAI211HDV2 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(B_inv, B );
	and SMC_I2(ZN_row1, A1_inv, B_inv );
	not SMC_I3(A2_inv, A2 );
	and SMC_I4(ZN_row2, A2_inv, B_inv );
	not SMC_I5(C_inv, C );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2, C_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOAI211HDV4 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(B_inv, B );
	and SMC_I2(ZN_row1, A1_inv, B_inv );
	not SMC_I3(A2_inv, A2 );
	and SMC_I4(ZN_row2, A2_inv, B_inv );
	not SMC_I5(C_inv, C );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2, C_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOAI211HDV8 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(B_inv, B );
	and SMC_I2(ZN_row1, A1_inv, B_inv );
	not SMC_I3(A2_inv, A2 );
	and SMC_I4(ZN_row2, A2_inv, B_inv );
	not SMC_I5(C_inv, C );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2, C_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOAI211HDVL ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(B_inv, B );
	and SMC_I2(ZN_row1, A1_inv, B_inv );
	not SMC_I3(A2_inv, A2 );
	and SMC_I4(ZN_row2, A2_inv, B_inv );
	not SMC_I5(C_inv, C );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2, C_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211HDV0 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A1, A2 );
  nor I1(ZN_temp, B, C, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211HDV1 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A1, A2 );
  nor I1(ZN_temp, B, C, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211HDV2 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A1, A2 );
  nor I1(ZN_temp, B, C, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211HDV4 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A1, A2 );
  nor I1(ZN_temp, B, C, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211HDV8 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A1, A2 );
  nor I1(ZN_temp, B, C, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI211HDVL ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A1, A2 );
  nor I1(ZN_temp, B, C, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21BHDV0 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, B1, B2 );
    not SMC_I1(OUT1, A );
    nor	SMC_I2(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(B1===1'b0 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21BHDV1 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, B1, B2 );
    not SMC_I1(OUT1, A );
    nor	SMC_I2(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(B1===1'b0 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21BHDV2 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, B1, B2 );
    not SMC_I1(OUT1, A );
    nor	SMC_I2(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(B1===1'b0 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21BHDV4 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, B1, B2 );
    not SMC_I1(OUT1, A );
    nor	SMC_I2(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(B1===1'b0 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21BHDV8 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, B1, B2 );
    not SMC_I1(OUT1, A );
    nor	SMC_I2(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(B1===1'b0 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21BHDVL ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, B1, B2 );
    not SMC_I1(OUT1, A );
    nor	SMC_I2(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(B1===1'b0 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21HDV0 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, A1, A2 );
    nor SMC_I1(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21HDV1 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, A1, A2 );
    nor SMC_I1(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21HDV12 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, A1, A2 );
    nor SMC_I1(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21HDV2 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, A1, A2 );
    nor SMC_I1(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21HDV4 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, A1, A2 );
    nor SMC_I1(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21HDV8 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, A1, A2 );
    nor SMC_I1(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI21HDVL ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    and SMC_I0(OUT0, A1, A2 );
    nor SMC_I1(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221HDV0 ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A2, A1 );
  and I1(out1, B2, B1 );
  nor I2(ZN_temp, C, out1, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221HDV1 ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A2, A1 );
  and I1(out1, B2, B1 );
  nor I2(ZN_temp, C, out1, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221HDV2 ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A2, A1 );
  and I1(out1, B2, B1 );
  nor I2(ZN_temp, C, out1, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221HDV4 ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A2, A1 );
  and I1(out1, B2, B1 );
  nor I2(ZN_temp, C, out1, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI221HDVL ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(out0, A2, A1 );
  and I1(out1, B2, B1 );
  nor I2(ZN_temp, C, out1, out0 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222HDV0 ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  and I2(outC, C2, C1 );
  nor I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222HDV1 ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  and I2(outC, C2, C1 );
  nor I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222HDV2 ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  and I2(outC, C2, C1 );
  nor I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222HDV4 ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  and I2(outC, C2, C1 );
  nor I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI222HDVL ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  and I2(outC, C2, C1 );
  nor I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI22HDV0 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI22HDV1 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI22HDV2 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI22HDV4 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI22HDV8 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI22HDVL ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A2, A1 );
  and I1(outB, B2, B1 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI31HDV0 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  nor I1(ZN_temp, B, outA );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI31HDV1 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  nor I1(ZN_temp, B, outA );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI31HDV2 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  nor I1(ZN_temp, B, outA );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI31HDV4 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  nor I1(ZN_temp, B, outA );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI31HDV8 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  nor I1(ZN_temp, B, outA );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI31HDVL ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  nor I1(ZN_temp, B, outA );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI32HDV0 ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI32HDV1 ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI32HDV2 ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI32HDV4 ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI32HDVL ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI33HDV0 ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2, B3 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI33HDV1 ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2, B3 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI33HDV2 ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2, B3 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI33HDV4 ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2, B3 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module AOI33HDVL ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  and I0(outA, A1, A2, A3 );
  and I1(outB, B1, B2, B3 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV0 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV0RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV1 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV12 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV12RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV16 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV16RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV1RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV2 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV20 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV20RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV24 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV24RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV2RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV3 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV32 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV32RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV3RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV4 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV4RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV6 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV6RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV8 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDV8RD ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module BUFHDVL ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKAND2HDV0 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKAND2HDV1 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKAND2HDV12 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKAND2HDV2 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKAND2HDV4 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKAND2HDV8 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    and SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV0 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV1 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV12 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV16 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV2 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV20 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV24 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV3 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV32 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV4 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV6 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKBUFHDV8 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV0 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV1 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV12 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV16 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV2 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV20 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV24 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV3 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV4 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV6 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKINHDV8 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not SMC_I0 (ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc I --> ZN
	 (I => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDV0 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDV1 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDV12 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDV16 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDV2 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDV3 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDV4 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDV8 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKNAND2HDVL ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand SMC_I0 (ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKXOR2HDV0 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKXOR2HDV1 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKXOR2HDV2 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKXOR2HDV4 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor SMC_I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL1HDV0 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL1HDV1 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL1HDV2 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL1HDV4 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL2HDV0 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL2HDV1 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL2HDV2 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL2HDV4 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL3HDV0 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL3HDV1 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL3HDV2 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL3HDV4 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL4HDV0 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL4HDV1 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL4HDV2 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DEL4HDV4 ( Z, I, VDD, VSS); 
input I;
inout VDD, VSS;
output Z;
wire Z_temp;

	buf SMC_I0(Z_temp, I );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc I --> Z
	 (I => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module F_DIODEHD2 ( A, VDD, VSS); 
input A;
inout VDD, VSS;


   `ifdef functional  //  functional //

   `else




   specify

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module F_DIODEHD4 ( A, VDD, VSS); 
input A;
inout VDD, VSS;


   `ifdef functional  //  functional //

   `else




   specify

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module F_DIODEHD8 ( A, VDD, VSS); 
input A;
inout VDD, VSS;


   `ifdef functional  //  functional //

   `else




   specify

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NAND4HDV0 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nand (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NAND4HDV1 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nand (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NAND4HDV2 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nand (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NAND4HDV4 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nand (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NAND4HDVL ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nand (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NOR4HDV0 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nor (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NOR4HDV1 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nor (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NOR4HDV2 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nor (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NOR4HDV4 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nor (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module I2NOR4HDVL ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not (A1x, A1 );
  not (A2x, A2 );
  nor (ZN_temp, A1x, A2x, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO21HDV0 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(B_bar, B );
    and I1(OUT0, A2, B_bar );
    and I2(OUT1, A1, B_bar );
    or  I3(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO21HDV1 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(B_bar, B );
    and I1(OUT0, A2, B_bar );
    and I2(OUT1, A1, B_bar );
    or  I3(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO21HDV2 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(B_bar, B );
    and I1(OUT0, A2, B_bar );
    and I2(OUT1, A1, B_bar );
    or  I3(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO21HDV4 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(B_bar, B );
    and I1(OUT0, A2, B_bar );
    and I2(OUT1, A1, B_bar );
    or  I3(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO21HDV8 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(B_bar, B );
    and I1(OUT0, A2, B_bar );
    and I2(OUT1, A1, B_bar );
    or  I3(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO21HDVL ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(B_bar, B );
    and I1(OUT0, A2, B_bar );
    and I2(OUT1, A1, B_bar );
    or  I3(ZN_temp, OUT0, OUT1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO22HDV0 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nor I0 (outA, A1, A2 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO22HDV1 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nor I0 (outA, A1, A2 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO22HDV2 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nor I0 (outA, A1, A2 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO22HDV4 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nor I0 (outA, A1, A2 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IAO22HDVL ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nor I0 (outA, A1, A2 );
  and I1(outB, B1, B2 );
  nor I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND2HDV0 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(A1_bar, A1 );
    nand I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND2HDV1 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(A1_bar, A1 );
    nand I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND2HDV12 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(A1_bar, A1 );
    nand I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND2HDV2 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(A1_bar, A1 );
    nand I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND2HDV4 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(A1_bar, A1 );
    nand I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND2HDV8 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(A1_bar, A1 );
    nand I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND2HDVL ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(A1_bar, A1 );
    nand I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND3HDV0 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND3HDV1 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND3HDV2 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND3HDV4 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND3HDV8 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND3HDVL ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND4HDV0 ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND4HDV1 ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND4HDV2 ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND4HDV4 ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INAND4HDVL ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nand I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV0 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV1 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV12 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV16 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV2 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV20 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV24 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV3 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV32 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV4 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV6 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDV8 ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INHDVL ( ZN, I, VDD, VSS); 
input I;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    not I0(ZN_temp, I );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> ZN 
	 (I => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR2HDV0 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not I0(A1_bar, A1 );
  nor I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR2HDV1 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not I0(A1_bar, A1 );
  nor I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR2HDV12 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not I0(A1_bar, A1 );
  nor I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR2HDV2 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not I0(A1_bar, A1 );
  nor I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR2HDV4 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not I0(A1_bar, A1 );
  nor I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR2HDV8 ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not I0(A1_bar, A1 );
  nor I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR2HDVL ( ZN, A1, B1, VDD, VSS); 
input A1, B1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  not I0(A1_bar, A1 );
  nor I1(ZN_temp, A1_bar, B1 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR3HDV0 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR3HDV1 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR3HDV2 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR3HDV4 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR3HDV8 ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR3HDVL ( ZN, A1, B1, B2, VDD, VSS); 
input A1, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR4HDV0 ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR4HDV1 ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR4HDV2 ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR4HDV4 ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module INOR4HDVL ( ZN, A1, B1, B2, B3, VDD, VSS); 
input A1, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not I0(A1_bar, A1 );
   nor I1(ZN_temp, A1_bar, B1, B2, B3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA21HDV0 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nand I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA21HDV1 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nand I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA21HDV2 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nand I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA21HDV4 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nand I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA21HDV8 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nand I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA21HDVL ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  nand I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA22HDV0 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA22HDV1 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA22HDV2 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA22HDV4 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module IOA22HDVL ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAJ23HDV0 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

	and SMC_I0(Z_row1, A1, A2 );
	and SMC_I1(Z_row2, A1, A3 );
	and SMC_I2(Z_row3, A2, A3 );
	or SMC_I3(Z_temp, Z_row1, Z_row2, Z_row3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	if(A2===1'b0 && A3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A2===1'b1 && A3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAJ23HDV1 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

	and SMC_I0(Z_row1, A1, A2 );
	and SMC_I1(Z_row2, A1, A3 );
	and SMC_I2(Z_row3, A2, A3 );
	or SMC_I3(Z_temp, Z_row1, Z_row2, Z_row3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	if(A2===1'b0 && A3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A2===1'b1 && A3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAJ23HDV2 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

	and SMC_I0(Z_row1, A1, A2 );
	and SMC_I1(Z_row2, A1, A3 );
	and SMC_I2(Z_row3, A2, A3 );
	or SMC_I3(Z_temp, Z_row1, Z_row2, Z_row3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	if(A2===1'b0 && A3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A2===1'b1 && A3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAJ23HDV4 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

	and SMC_I0(Z_row1, A1, A2 );
	and SMC_I1(Z_row2, A1, A3 );
	and SMC_I2(Z_row3, A2, A3 );
	or SMC_I3(Z_temp, Z_row1, Z_row2, Z_row3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	if(A2===1'b0 && A3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A2===1'b1 && A3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAJ23HDV8 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

	and SMC_I0(Z_row1, A1, A2 );
	and SMC_I1(Z_row2, A1, A3 );
	and SMC_I2(Z_row3, A2, A3 );
	or SMC_I3(Z_temp, Z_row1, Z_row2, Z_row3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	if(A2===1'b0 && A3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A2===1'b1 && A3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAJ23HDVL ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

	and SMC_I0(Z_row1, A1, A2 );
	and SMC_I1(Z_row2, A1, A3 );
	and SMC_I2(Z_row3, A2, A3 );
	or SMC_I3(Z_temp, Z_row1, Z_row2, Z_row3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	if(A2===1'b0 && A3===1'b1)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A2===1'b1 && A3===1'b0)
	// arc A1 --> Z
	 (A1 => Z) = (1.0,1.0);

	if(A1===1'b0 && A3===1'b1)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b1 && A3===1'b0)
	// arc A2 --> Z
	 (A2 => Z) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc A3 --> Z
	 (A3 => Z) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAOI222HDV0 ( ZN, A, B, C, VDD, VSS); 
input A, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   and I0(outAB, A, B );
   and I1(outBC, B, C );
   and I2(outAC, A, C );
   nor I3(ZN_temp, outAB, outBC, outAC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && C===1'b1) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(B===1'b1 && C===1'b0) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && C===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && C===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAOI222HDV1 ( ZN, A, B, C, VDD, VSS); 
input A, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   and I0(outAB, A, B );
   and I1(outBC, B, C );
   and I2(outAC, A, C );
   nor I3(ZN_temp, outAB, outBC, outAC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && C===1'b1) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(B===1'b1 && C===1'b0) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && C===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && C===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAOI222HDV2 ( ZN, A, B, C, VDD, VSS); 
input A, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   and I0(outAB, A, B );
   and I1(outBC, B, C );
   and I2(outAC, A, C );
   nor I3(ZN_temp, outAB, outBC, outAC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && C===1'b1) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(B===1'b1 && C===1'b0) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && C===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && C===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAOI222HDV4 ( ZN, A, B, C, VDD, VSS); 
input A, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   and I0(outAB, A, B );
   and I1(outBC, B, C );
   and I2(outAC, A, C );
   nor I3(ZN_temp, outAB, outBC, outAC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && C===1'b1) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(B===1'b1 && C===1'b0) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && C===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && C===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MAOI222HDVL ( ZN, A, B, C, VDD, VSS); 
input A, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   and I0(outAB, A, B );
   and I1(outBC, B, C );
   and I2(outAC, A, C );
   nor I3(ZN_temp, outAB, outBC, outAC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B===1'b0 && C===1'b1) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(B===1'b1 && C===1'b0) 
	// arc A --> ZN 
	 (A => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && C===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && C===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A===1'b0 && B===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A===1'b1 && B===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV0 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV1 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV12 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV16 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV2 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV24 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV3 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV4 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDV8 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND2HDVL ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nand I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3BBHDV0 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      not  I1(A1_inv, A1 );
      not  I2(A2_inv, A2 );
      and  I3(OUT0, A1_inv, A2_inv );
      nand I0(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3BBHDV1 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      not  I1(A1_inv, A1 );
      not  I2(A2_inv, A2 );
      and  I3(OUT0, A1_inv, A2_inv );
      nand I0(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3BBHDV2 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      not  I1(A1_inv, A1 );
      not  I2(A2_inv, A2 );
      and  I3(OUT0, A1_inv, A2_inv );
      nand I0(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3BBHDV4 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      not  I1(A1_inv, A1 );
      not  I2(A2_inv, A2 );
      and  I3(OUT0, A1_inv, A2_inv );
      nand I0(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3BBHDV8 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      not  I1(A1_inv, A1 );
      not  I2(A2_inv, A2 );
      and  I3(OUT0, A1_inv, A2_inv );
      nand I0(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3BBHDVL ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      not  I1(A1_inv, A1 );
      not  I2(A2_inv, A2 );
      and  I3(OUT0, A1_inv, A2_inv );
      nand I0(ZN_temp, OUT0, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3HDV0 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      nand I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3HDV1 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      nand I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3HDV12 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      nand I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3HDV2 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      nand I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3HDV3 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      nand I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3HDV4 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      nand I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3HDV8 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      nand I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND3HDVL ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

      nand I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND4HDV0 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND4HDV1 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND4HDV2 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND4HDV3 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND4HDV4 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND4HDV8 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NAND4HDVL ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nand I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDV0 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDV1 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDV12 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDV16 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDV2 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDV3 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDV4 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDV8 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR2HDVL ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    nor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3BBHDV0 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not  I1(A1_inv, A1 );
   not  I2(A2_inv, A2 );
   nor  I0(ZN_temp, A1_inv, A2_inv, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
  	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3BBHDV1 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not  I1(A1_inv, A1 );
   not  I2(A2_inv, A2 );
   nor  I0(ZN_temp, A1_inv, A2_inv, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
  	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3BBHDV2 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not  I1(A1_inv, A1 );
   not  I2(A2_inv, A2 );
   nor  I0(ZN_temp, A1_inv, A2_inv, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
  	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3BBHDV4 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not  I1(A1_inv, A1 );
   not  I2(A2_inv, A2 );
   nor  I0(ZN_temp, A1_inv, A2_inv, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
  	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3BBHDV8 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not  I1(A1_inv, A1 );
   not  I2(A2_inv, A2 );
   nor  I0(ZN_temp, A1_inv, A2_inv, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
  	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3BBHDVL ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   not  I1(A1_inv, A1 );
   not  I2(A2_inv, A2 );
   nor  I0(ZN_temp, A1_inv, A2_inv, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
  	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3HDV0 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor  I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3HDV1 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor  I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3HDV12 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor  I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3HDV2 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor  I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3HDV3 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor  I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3HDV4 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor  I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3HDV8 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor  I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR3HDVL ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor  I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR4HDV0 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR4HDV1 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR4HDV2 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR4HDV3 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR4HDV4 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR4HDV8 ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NOR4HDVL ( ZN, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   nor I0(ZN_temp, A1, A2, A3, A4 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	// arc A4 --> ZN 
	 (A4 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA211HDV0 ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or   I0(outA, A1, A2 );
   and  I1(Z_temp, B, C, outA );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA211HDV1 ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or   I0(outA, A1, A2 );
   and  I1(Z_temp, B, C, outA );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA211HDV2 ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or   I0(outA, A1, A2 );
   and  I1(Z_temp, B, C, outA );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA211HDV4 ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or   I0(outA, A1, A2 );
   and  I1(Z_temp, B, C, outA );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA211HDVL ( Z, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or   I0(outA, A1, A2 );
   and  I1(Z_temp, B, C, outA );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA21HDV0 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA21HDV1 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA21HDV2 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA21HDV4 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA21HDV8 ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA21HDVL ( Z, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA221HDV0 ( Z, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   and I2(Z_temp, outA, outB, C );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA221HDV1 ( Z, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   and I2(Z_temp, outA, outB, C );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA221HDV2 ( Z, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   and I2(Z_temp, outA, outB, C );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA221HDV4 ( Z, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output Z;
wire Z_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   and I2(Z_temp, outA, outB, C );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> Z 
	 (C => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA222HDV0 ( Z, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output Z;
wire Z_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   or  I2(outC, C1, C2 );
   and I3(Z_temp, outA, outB, outC );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA222HDV1 ( Z, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output Z;
wire Z_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   or  I2(outC, C1, C2 );
   and I3(Z_temp, outA, outB, outC );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA222HDV2 ( Z, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output Z;
wire Z_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   or  I2(outC, C1, C2 );
   and I3(Z_temp, outA, outB, outC );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA222HDV4 ( Z, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output Z;
wire Z_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   or  I2(outC, C1, C2 );
   and I3(Z_temp, outA, outB, outC );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> Z 
	 (C1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> Z 
	 (C2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA22HDV0 ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA22HDV1 ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA22HDV2 ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA22HDV4 ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA22HDVL ( Z, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA31HDV0 ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA31HDV1 ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA31HDV2 ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA31HDV4 ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA31HDVL ( Z, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    and I1(Z_temp, outA, B );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> Z 
	 (B => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA32HDV0 ( Z, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2, A3 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA32HDV1 ( Z, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2, A3 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA32HDV2 ( Z, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2, A3 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA32HDV4 ( Z, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output Z;
wire Z_temp;

  or  I0(outA, A1, A2, A3 );
  or  I1(outB, B1, B2 );
  and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA33HDV0 ( Z, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    or  I1(outB, B1, B2, B3 );
    and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA33HDV1 ( Z, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    or  I1(outB, B1, B2, B3 );
    and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA33HDV2 ( Z, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    or  I1(outB, B1, B2, B3 );
    and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OA33HDV4 ( Z, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or  I0(outA, A1, A2, A3 );
    or  I1(outB, B1, B2, B3 );
    and I2(Z_temp, outA, outB );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> Z 
	 (B1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> Z 
	 (B2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> Z 
	 (B3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI211HDV0 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI211HDV1 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI211HDV2 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI211HDV4 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI211HDV8 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI211HDVL ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21BHDV0 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outB, B1, B2 );
  not  I2(A_inv, A );
  nand I1(ZN_temp, outB, A_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21BHDV1 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outB, B1, B2 );
  not  I2(A_inv, A );
  nand I1(ZN_temp, outB, A_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21BHDV2 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outB, B1, B2 );
  not  I2(A_inv, A );
  nand I1(ZN_temp, outB, A_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21BHDV4 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outB, B1, B2 );
  not  I2(A_inv, A );
  nand I1(ZN_temp, outB, A_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21BHDV8 ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outB, B1, B2 );
  not  I2(A_inv, A );
  nand I1(ZN_temp, outB, A_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21BHDVL ( ZN, A, B1, B2, VDD, VSS); 
input A, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outB, B1, B2 );
  not  I2(A_inv, A );
  nand I1(ZN_temp, outB, A_inv );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 	if(B1===1'b0 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b0)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	if(B1===1'b1 && B2===1'b1)
	// arc A --> ZN
	 (A => ZN) = (1.0,1.0);

	// arc B1 --> ZN
	 (B1 => ZN) = (1.0,1.0);

	// arc B2 --> ZN
	 (B2 => ZN) = (1.0,1.0);
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21HDV0 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21HDV1 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21HDV12 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21HDV16 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21HDV2 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21HDV4 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21HDV8 ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI21HDVL ( ZN, A1, A2, B, VDD, VSS); 
input A1, A2, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  or   I0(outA, A1, A2 );
  nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221HDV0 ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221HDV1 ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221HDV2 ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221HDV4 ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI221HDVL ( ZN, A1, A2, B1, B2, C, VDD, VSS); 
input A1, A2, B1, B2, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or  I0(outA, A1, A2 );
   or  I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB, C );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C --> ZN 
	 (C => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222HDV0 ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   or   I2(outC, C1, C2 );
   nand I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222HDV1 ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   or   I2(outC, C1, C2 );
   nand I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222HDV2 ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   or   I2(outC, C1, C2 );
   nand I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222HDV4 ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   or   I2(outC, C1, C2 );
   nand I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI222HDVL ( ZN, A1, A2, B1, B2, C1, C2, VDD, VSS); 
input A1, A2, B1, B2, C1, C2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   or   I2(outC, C1, C2 );
   nand I3(ZN_temp, outA, outB, outC );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b0 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && C1===1'b1 && C2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C1 --> ZN 
	 (C1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1) 
	// arc C2 --> ZN 
	 (C2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22HDV0 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22HDV1 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22HDV2 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22HDV4 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22HDV8 ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI22HDVL ( ZN, A1, A2, B1, B2, VDD, VSS); 
input A1, A2, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31HDV0 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31HDV1 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31HDV2 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31HDV4 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31HDV8 ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI31HDVL ( ZN, A1, A2, A3, B, VDD, VSS); 
input A1, A2, A3, B;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   nand I1(ZN_temp, outA, B );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B --> ZN 
	 (B => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32HDV0 ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32HDV1 ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32HDV2 ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32HDV4 ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI32HDVL ( ZN, A1, A2, A3, B1, B2, VDD, VSS); 
input A1, A2, A3, B1, B2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33HDV0 ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2, B3 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33HDV1 ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2, B3 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33HDV2 ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2, B3 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33HDV4 ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2, B3 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAI33HDVL ( ZN, A1, A2, A3, B1, B2, B3, VDD, VSS); 
input A1, A2, A3, B1, B2, B3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   or   I0(outA, A1, A2, A3 );
   or   I1(outB, B1, B2, B3 );
   nand I2(ZN_temp, outA, outB );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b0 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b0 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(B1===1'b1 && B2===1'b1 && B3===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B1 --> ZN 
	 (B1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B2 --> ZN 
	 (B2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b0) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1 && A3===1'b1) 
	// arc B3 --> ZN 
	 (B3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAOI211HDV0 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(A2_inv, A2 );
	not SMC_I2(C_inv, C );
	and SMC_I3(ZN_row1, A1_inv, A2_inv, C_inv );
	not SMC_I4(B_inv, B );
	and SMC_I5(ZN_row2, B_inv, C_inv );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAOI211HDV1 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(A2_inv, A2 );
	not SMC_I2(C_inv, C );
	and SMC_I3(ZN_row1, A1_inv, A2_inv, C_inv );
	not SMC_I4(B_inv, B );
	and SMC_I5(ZN_row2, B_inv, C_inv );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAOI211HDV2 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(A2_inv, A2 );
	not SMC_I2(C_inv, C );
	and SMC_I3(ZN_row1, A1_inv, A2_inv, C_inv );
	not SMC_I4(B_inv, B );
	and SMC_I5(ZN_row2, B_inv, C_inv );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAOI211HDV4 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(A2_inv, A2 );
	not SMC_I2(C_inv, C );
	and SMC_I3(ZN_row1, A1_inv, A2_inv, C_inv );
	not SMC_I4(B_inv, B );
	and SMC_I5(ZN_row2, B_inv, C_inv );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAOI211HDV8 ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(A2_inv, A2 );
	not SMC_I2(C_inv, C );
	and SMC_I3(ZN_row1, A1_inv, A2_inv, C_inv );
	not SMC_I4(B_inv, B );
	and SMC_I5(ZN_row2, B_inv, C_inv );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OAOI211HDVL ( ZN, A1, A2, B, C, VDD, VSS); 
input A1, A2, B, C;
inout VDD, VSS;
output ZN;
wire ZN_temp;

	not SMC_I0(A1_inv, A1 );
	not SMC_I1(A2_inv, A2 );
	not SMC_I2(C_inv, C );
	and SMC_I3(ZN_row1, A1_inv, A2_inv, C_inv );
	not SMC_I4(B_inv, B );
	and SMC_I5(ZN_row2, B_inv, C_inv );
	or SMC_I6(ZN_temp, ZN_row1, ZN_row2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

	// arc A1 --> ZN
	 (A1 => ZN) = (1.0,1.0);

	// arc A2 --> ZN
	 (A2 => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1)
	// arc B --> ZN
	 (B => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b0 && B===1'b1)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b0 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b0 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

	if(A1===1'b1 && A2===1'b1 && B===1'b0)
	// arc C --> ZN
	 (C => ZN) = (1.0,1.0);

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV0 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV0RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV1 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV12 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV12RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV16 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV16RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV1RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV2 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV2RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV4 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV4RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV8 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDV8RD ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR2HDVL ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV0 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV0RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV1 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV1RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV2 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV2RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV4 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV4RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV8 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDV8RD ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR3HDVL ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

    or (Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR4HDV0 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(OUT0, A4 );
    buf I1(OUT1, A2 );
    buf I2(OUT2, A3 );
    buf I3(OUT3, A1 );
    or  I4(Z_temp, OUT0, OUT1, OUT2, OUT3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR4HDV1 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(OUT0, A4 );
    buf I1(OUT1, A2 );
    buf I2(OUT2, A3 );
    buf I3(OUT3, A1 );
    or  I4(Z_temp, OUT0, OUT1, OUT2, OUT3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR4HDV2 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(OUT0, A4 );
    buf I1(OUT1, A2 );
    buf I2(OUT2, A3 );
    buf I3(OUT3, A1 );
    or  I4(Z_temp, OUT0, OUT1, OUT2, OUT3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR4HDV4 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(OUT0, A4 );
    buf I1(OUT1, A2 );
    buf I2(OUT2, A3 );
    buf I3(OUT3, A1 );
    or  I4(Z_temp, OUT0, OUT1, OUT2, OUT3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR4HDV8 ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(OUT0, A4 );
    buf I1(OUT1, A2 );
    buf I2(OUT2, A3 );
    buf I3(OUT3, A1 );
    or  I4(Z_temp, OUT0, OUT1, OUT2, OUT3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module OR4HDVL ( Z, A1, A2, A3, A4, VDD, VSS); 
input A1, A2, A3, A4;
inout VDD, VSS;
output Z;
wire Z_temp;

    buf I0(OUT0, A4 );
    buf I1(OUT1, A2 );
    buf I2(OUT2, A3 );
    buf I3(OUT3, A1 );
    or  I4(Z_temp, OUT0, OUT1, OUT2, OUT3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	// arc A4 --> Z 
	 (A4 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module PULLHD0 ( Z, VDD, VSS); 
inout VDD, VSS;
output Z;
wire Z_temp;

	assign Z = 1'b0; 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module PULLHD1 ( Z, VDD, VSS); 
inout VDD, VSS;
output Z;
wire Z_temp;

	assign Z = 1'b1; 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
   `ifdef functional  //  functional //

   `else




   specify

   endspecify

  `endif // functional //

endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV0 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV1 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV12 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV16 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV2 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV20 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV24 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV3 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV4 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV6 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module TBUFHDV8 ( Z, I, OE, VDD, VSS); 
input I, OE;
inout VDD, VSS;
output Z;
wire Z_temp;

  bufif1 I0(Z_temp, I, OE );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc I --> Z 
	 (I => Z) = (1.0,1.0); 
 
	// arc OE --> Z 
	 (OE => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2CHDV0 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2CHDV1 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2CHDV2 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2CHDV4 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2CHDV8 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2CHDVL ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2HDV0 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2HDV1 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2HDV2 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2HDV4 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2HDV8 ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR2HDVL ( ZN, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output ZN;
wire ZN_temp;

    xnor I0(ZN_temp, A1, A2 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (ZN:A1) 
	 (posedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (ZN:A1) 
	 (negedge A1 => (ZN:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (ZN:A2) 
	 (posedge A2 => (ZN:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (ZN:A2) 
	 (negedge A2 => (ZN:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR3HDV0 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   xnor I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR3HDV1 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   xnor I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR3HDV2 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   xnor I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR3HDV4 ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   xnor I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XNOR3HDVL ( ZN, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   xnor I0(ZN_temp, A1, A2, A3 );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> ZN 
	 (A1 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> ZN 
	 (A2 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> ZN 
	 (A3 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2CHDV0 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2CHDV1 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2CHDV2 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2CHDV4 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2CHDV8 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2CHDVL ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2HDV0 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2HDV1 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2HDV2 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2HDV4 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2HDV8 ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR2HDVL ( Z, A1, A2, VDD, VSS); 
input A1, A2;
inout VDD, VSS;
output Z;
wire Z_temp;

    xor I0(Z_temp, A1, A2 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc posedge A1 --> (Z:A1) 
	 (posedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc negedge A1 --> (Z:A1) 
	 (negedge A1 => (Z:A1)) = (1.0,1.0); 
 
	// arc posedge A2 --> (Z:A2) 
	 (posedge A2 => (Z:A2)) = (1.0,1.0); 
 
	// arc negedge A2 --> (Z:A2) 
	 (negedge A2 => (Z:A2)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3HDV0 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

   xor I0(Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3HDV1 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

   xor I0(Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3HDV2 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

   xor I0(Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3HDV4 ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

   xor I0(Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module XOR3HDVL ( Z, A1, A2, A3, VDD, VSS); 
input A1, A2, A3;
inout VDD, VSS;
output Z;
wire Z_temp;

   xor I0(Z_temp, A1, A2, A3 );
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(A2===1'b0 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b0 && A3===1'b0) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A2===1'b1 && A3===1'b1) 
	// arc A1 --> Z 
	 (A1 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A3===1'b0) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A3===1'b1) 
	// arc A2 --> Z 
	 (A2 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b0 && A2===1'b0) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
	if(A1===1'b1 && A2===1'b1) 
	// arc A3 --> Z 
	 (A3 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHAQHDV0 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE; 
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  udp_tlat_PWR I4 (n1, xE, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I5 (cond0, n1 );
  not      I6 (nTE, TE );
  and      I7 (n0, nTE, cond0 );
  or       I8 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHAQHDV1 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE; 
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  udp_tlat_PWR I4 (n1, xE, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I5 (cond0, n1 );
  not      I6 (nTE, TE );
  and      I7 (n0, nTE, cond0 );
  or       I8 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHAQHDV2 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE; 
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  udp_tlat_PWR I4 (n1, xE, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I5 (cond0, n1 );
  not      I6 (nTE, TE );
  and      I7 (n0, nTE, cond0 );
  or       I8 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHAQHDV4 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE; 
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  udp_tlat_PWR I4 (n1, xE, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I5 (cond0, n1 );
  not      I6 (nTE, TE );
  and      I7 (n0, nTE, cond0 );
  or       I8 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHAQHDV8 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE; 
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  udp_tlat_PWR I4 (n1, xE, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I5 (cond0, n1 );
  not      I6 (nTE, TE );
  and      I7 (n0, nTE, cond0 );
  or       I8 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHQHDV0 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  or       I4 (n0, xE, xTE );
  udp_tlat_PWR I5 (n1, n0, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I6 (cond0, n1 );
  or       I7 (Q_temp, cond0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
  endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHQHDV1 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  or       I4 (n0, xE, xTE );
  udp_tlat_PWR I5 (n1, n0, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I6 (cond0, n1 );
  or       I7 (Q_temp, cond0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
  endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHQHDV2 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  or       I4 (n0, xE, xTE );
  udp_tlat_PWR I5 (n1, n0, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I6 (cond0, n1 );
  or       I7 (Q_temp, cond0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
  endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHQHDV4 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  or       I4 (n0, xE, xTE );
  udp_tlat_PWR I5 (n1, n0, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I6 (cond0, n1 );
  or       I7 (Q_temp, cond0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
  endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLAHQHDV8 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  not      I3 (nclk, dCK );
  or       I4 (n0, xE, xTE );
  udp_tlat_PWR I5 (n1, n0, nclk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not      I6 (cond0, n1 );
  or       I7 (Q_temp, cond0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(negedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
  endspecify 
 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANAQHDV0 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, TE );
  buf      I2 (xE, dE );
  udp_tlat_PWR I3 (n1, xE, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  or       I4 (n0, n1, xTE );
  and      I5 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANAQHDV1 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, TE );
  buf      I2 (xE, dE );
  udp_tlat_PWR I3 (n1, xE, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  or       I4 (n0, n1, xTE );
  and      I5 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANAQHDV2 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, TE );
  buf      I2 (xE, dE );
  udp_tlat_PWR I3 (n1, xE, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  or       I4 (n0, n1, xTE );
  and      I5 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANAQHDV4 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, TE );
  buf      I2 (xE, dE );
  udp_tlat_PWR I3 (n1, xE, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  or       I4 (n0, n1, xTE );
  and      I5 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANAQHDV8 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, TE );
  buf      I2 (xE, dE );
  udp_tlat_PWR I3 (n1, xE, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  or       I4 (n0, n1, xTE );
  and      I5 (Q_temp, n0, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&&(ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
   endspecify 
  `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV0 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV1 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV12 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV16 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV2 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV20 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV24 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV3 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV4 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV6 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKLANQHDV8 ( Q, CK, E, TE, VDD, VSS); 
input CK, E, TE;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
wire ENABLE_NOT_TE;
wire ENABLE_NOT_E;
assign ENABLE_NOT_TE = (!TE) ? 1'b1:1'b0;
assign ENABLE_NOT_E = (!E) ? 1'b1:1'b0;
  buf      I0 (clk, dCK );
  buf      I1 (xTE, dTE );
  buf      I2 (xE, dE );
  or       I3 (n0, xE, xTE );
  udp_tlat_PWR I4 (n1, n0, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  and      I5 (Q_temp, n1, clk );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
 
   specify 
 
 
 	if(E===1'b0 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 

	if(E===1'b0 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b0) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0); 
 
	if(E===1'b1 && TE===1'b1) 
	// arc CK --> Q 
	 (CK => Q) = (1.0,1.0);
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_TE === 1'b1), posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), negedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_E === 1'b1), posedge TE, 1.0, 1.0, NOTIFIER, , , dCK, dTE); 
 
 
 
 
        endspecify 
       `endif 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKMUX2HDV0 ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKMUX2HDV1 ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKMUX2HDV2 ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module CLKMUX2HDV4 ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DGRNQHDV0 ( Q, CK, D, RN, VDD, VSS); 
input CK, D, RN;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN, EN; 
  buf       X0 (xRN, dRN );
  buf       IC (clk, dCK );
  udp_edfft_PWR I0 (n0, dD, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER ); 
  buf       I1 (Q_temp, n0 );
  and       I4 (Deff, dD, xRN );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
        $setuphold(posedge CK, posedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DGRNQHDV2 ( Q, CK, D, RN, VDD, VSS); 
input CK, D, RN;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN, EN; 
  buf       X0 (xRN, dRN );
  buf       IC (clk, dCK );
  udp_edfft_PWR I0 (n0, dD, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER ); 
  buf       I1 (Q_temp, n0 );
  and       I4 (Deff, dD, xRN );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
        $setuphold(posedge CK, posedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DGRNQHDV4 ( Q, CK, D, RN, VDD, VSS); 
input CK, D, RN;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN, EN; 
  buf       X0 (xRN, dRN );
  buf       IC (clk, dCK );
  udp_edfft_PWR I0 (n0, dD, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER ); 
  buf       I1 (Q_temp, n0 );
  and       I4 (Deff, dD, xRN );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
        $setuphold(posedge CK, posedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DGRNQHDV8 ( Q, CK, D, RN, VDD, VSS); 
input CK, D, RN;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN, EN; 
  buf       X0 (xRN, dRN );
  buf       IC (clk, dCK );
  udp_edfft_PWR I0 (n0, dD, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER ); 
  buf       I1 (Q_temp, n0 );
  and       I4 (Deff, dD, xRN );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
        $setuphold(posedge CK, posedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DGRNQNHDV0 ( QN, CK, D, RN, VDD, VSS); 
input CK, D, RN;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN, EN; 
  buf       X0 (xRN, dRN );
  buf       IC (clk, dCK );
  udp_edfft_PWR I0 (n0, dD, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER ); 
  not       I2 (QN_temp, n0 );
  and       I4 (Deff, dD, xRN );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
        $setuphold(posedge CK, posedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DGRNQNHDV2 ( QN, CK, D, RN, VDD, VSS); 
input CK, D, RN;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN, EN; 
  buf       X0 (xRN, dRN );
  buf       IC (clk, dCK );
  udp_edfft_PWR I0 (n0, dD, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER ); 
  not       I2 (QN_temp, n0 );
  and       I4 (Deff, dD, xRN );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
        $setuphold(posedge CK, posedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DGRNQNHDV4 ( QN, CK, D, RN, VDD, VSS); 
input CK, D, RN;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN, EN; 
  buf       X0 (xRN, dRN );
  buf       IC (clk, dCK );
  udp_edfft_PWR I0 (n0, dD, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER ); 
  not       I2 (QN_temp, n0 );
  and       I4 (Deff, dD, xRN );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
        $setuphold(posedge CK, posedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DGRNQNHDV8 ( QN, CK, D, RN, VDD, VSS); 
input CK, D, RN;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN, EN; 
  buf       X0 (xRN, dRN );
  buf       IC (clk, dCK );
  udp_edfft_PWR I0 (n0, dD, clk, xRN, xSN, EN, VDD, VSS, NOTIFIER ); 
  not       I2 (QN_temp, n0 );
  and       I4 (Deff, dD, xRN );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
        $setuphold(posedge CK, posedge RN, 1.0, 1.0, NOTIFIER, , , dCK, dRN); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DQHDV0 ( Q, CK, D, VDD, VSS); 
input CK, D;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DQHDV2 ( Q, CK, D, VDD, VSS); 
input CK, D;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DQHDV4 ( Q, CK, D, VDD, VSS); 
input CK, D;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DQHDV8 ( Q, CK, D, VDD, VSS); 
input CK, D;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DQNHDV0 ( QN, CK, D, VDD, VSS); 
input CK, D;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DQNHDV2 ( QN, CK, D, VDD, VSS); 
input CK, D;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DQNHDV4 ( QN, CK, D, VDD, VSS); 
input CK, D;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DQNHDV8 ( QN, CK, D, VDD, VSS); 
input CK, D;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK, negedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
        $setuphold(posedge CK, posedge D, 1.0, 1.0, NOTIFIER, , , dCK, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRNQHDV0 (D, RDN, CK, Q, VDD, VSS); 
  input D, RDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRNQHDV2 (D, RDN, CK, Q, VDD, VSS); 
  input D, RDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRNQHDV4 (D, RDN, CK, Q, VDD, VSS); 
  input D, RDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRNQHDV8 (D, RDN, CK, Q, VDD, VSS); 
  input D, RDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRNQNHDV0 (D, RDN, CK, QN, VDD, VSS); 
  input D, RDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRNQNHDV2 (D, RDN, CK, QN, VDD, VSS); 
  input D, RDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRNQNHDV4 (D, RDN, CK, QN, VDD, VSS); 
  input D, RDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRNQNHDV8 (D, RDN, CK, QN, VDD, VSS); 
  input D, RDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRQHDV0 (D, RD, CK, Q, VDD, VSS); 
  input D, RD, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(ENABLE_NOT_RD,dRD);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), negedge RD &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRQHDV2 (D, RD, CK, Q, VDD, VSS); 
  input D, RD, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(ENABLE_NOT_RD,dRD);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), negedge RD &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRQHDV4 (D, RD, CK, Q, VDD, VSS); 
  input D, RD, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(ENABLE_NOT_RD,dRD);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), negedge RD &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRQHDV8 (D, RD, CK, Q, VDD, VSS); 
  input D, RD, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(ENABLE_NOT_RD,dRD);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), negedge RD &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRQNHDV0 (D, RD, CK, QN, VDD, VSS); 
  input D, RD, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(ENABLE_NOT_RD,dRD);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), negedge RD &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRQNHDV2 (D, RD, CK, QN, VDD, VSS); 
  input D, RD, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(ENABLE_NOT_RD,dRD);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), negedge RD &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRQNHDV4 (D, RD, CK, QN, VDD, VSS); 
  input D, RD, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(ENABLE_NOT_RD,dRD);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), negedge RD &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRQNHDV8 (D, RD, CK, QN, VDD, VSS); 
  input D, RD, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(ENABLE_NOT_RD,dRD);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge D &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D === 1'b1), negedge RD &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRSNQHDV0 (D, RDN, SDN, CK, Q, VDD, VSS); 
  input D, RDN, SDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRSNQHDV2 (D, RDN, SDN, CK, Q, VDD, VSS); 
  input D, RDN, SDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRSNQHDV4 (D, RDN, SDN, CK, Q, VDD, VSS); 
  input D, RDN, SDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRSNQHDV8 (D, RDN, SDN, CK, Q, VDD, VSS); 
  input D, RDN, SDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRSNQNHDV0 (D, RDN, SDN, CK, QN, VDD, VSS); 
  input D, RDN, SDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRSNQNHDV2 (D, RDN, SDN, CK, QN, VDD, VSS); 
  input D, RDN, SDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRSNQNHDV4 (D, RDN, SDN, CK, QN, VDD, VSS); 
  input D, RDN, SDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DRSNQNHDV8 (D, RDN, SDN, CK, QN, VDD, VSS); 
  input D, RDN, SDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DSNQHDV0 (D, SDN, CK, Q, VDD, VSS); 
  input D, SDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);


        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DSNQHDV2 (D, SDN, CK, Q, VDD, VSS); 
  input D, SDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);


        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DSNQHDV4 (D, SDN, CK, Q, VDD, VSS); 
  input D, SDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);


        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DSNQHDV8 (D, SDN, CK, Q, VDD, VSS); 
  input D, SDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);


        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DSNQNHDV0 (D, SDN, CK, QN, VDD, VSS); 
  input D, SDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DSNQNHDV2 (D, SDN, CK, QN, VDD, VSS); 
  input D, SDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DSNQNHDV4 (D, SDN, CK, QN, VDD, VSS); 
  input D, SDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DSNQNHDV8 (D, SDN, CK, QN, VDD, VSS); 
  input D, SDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DXHDV0 ( Q, QN, CK, DA, DB, SA, VDD, VSS); 
input CK, DA, DB, SA;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_mux2_PWR (d, dDB, dDA, dSA ,VDD, VSS); 
  udp_dff_PWR I0 (n0, d, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_SA,dSA); 
 
    not SMC_I7(ENABLE_NOT_SA,dSA); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : DA))  = (1.0,1.0); 
 
	// arc CK --> QN 
	(posedge CK => (QN : DA))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_SA === 1'b1), 
            negedge DA &&& (ENABLE_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
        $setuphold(posedge CK &&& (ENABLE_SA === 1'b1), 
            posedge DA &&& (ENABLE_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA === 1'b1), 
            negedge DB &&& (ENABLE_NOT_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA === 1'b1), 
            posedge DB &&& (ENABLE_NOT_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
 
 
        $setuphold(posedge CK, negedge SA, 1.0, 1.0, NOTIFIER, , , dCK, dSA); 
 
        $setuphold(posedge CK, posedge SA, 1.0, 1.0, NOTIFIER, , , dCK, dSA); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DXHDV2 ( Q, QN, CK, DA, DB, SA, VDD, VSS); 
input CK, DA, DB, SA;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_mux2_PWR (d, dDB, dDA, dSA ,VDD, VSS); 
  udp_dff_PWR I0 (n0, d, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_SA,dSA); 
 
    not SMC_I7(ENABLE_NOT_SA,dSA); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : DA))  = (1.0,1.0); 
 
	// arc CK --> QN 
	(posedge CK => (QN : DA))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_SA === 1'b1), 
            negedge DA &&& (ENABLE_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
        $setuphold(posedge CK &&& (ENABLE_SA === 1'b1), 
            posedge DA &&& (ENABLE_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA === 1'b1), 
            negedge DB &&& (ENABLE_NOT_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA === 1'b1), 
            posedge DB &&& (ENABLE_NOT_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
 
 
        $setuphold(posedge CK, negedge SA, 1.0, 1.0, NOTIFIER, , , dCK, dSA); 
 
        $setuphold(posedge CK, posedge SA, 1.0, 1.0, NOTIFIER, , , dCK, dSA); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module DXHDV4 ( Q, QN, CK, DA, DB, SA, VDD, VSS); 
input CK, DA, DB, SA;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  buf     IC (clk, dCK );
  udp_mux2_PWR (d, dDB, dDA, dSA ,VDD, VSS); 
  udp_dff_PWR I0 (n0, d, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_SA,dSA); 
 
    not SMC_I7(ENABLE_NOT_SA,dSA); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : DA))  = (1.0,1.0); 
 
	// arc CK --> QN 
	(posedge CK => (QN : DA))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_SA === 1'b1), 
            negedge DA &&& (ENABLE_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
        $setuphold(posedge CK &&& (ENABLE_SA === 1'b1), 
            posedge DA &&& (ENABLE_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA === 1'b1), 
            negedge DB &&& (ENABLE_NOT_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA === 1'b1), 
            posedge DB &&& (ENABLE_NOT_SA === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
 
 
        $setuphold(posedge CK, negedge SA, 1.0, 1.0, NOTIFIER, , , dCK, dSA); 
 
        $setuphold(posedge CK, posedge SA, 1.0, 1.0, NOTIFIER, , , dCK, dSA); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDQHDV0 ( Q, CK, D, E, VDD, VSS); 
input CK, D, E;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  buf     B1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_E,dE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            negedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            posedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK, posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDQHDV2 ( Q, CK, D, E, VDD, VSS); 
input CK, D, E;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  buf     B1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_E,dE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            negedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            posedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK, posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDQHDV4 ( Q, CK, D, E, VDD, VSS); 
input CK, D, E;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  buf     B1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_E,dE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            negedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            posedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK, posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDQHDV8 ( Q, CK, D, E, VDD, VSS); 
input CK, D, E;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  buf     B1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_E,dE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            negedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            posedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK, posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDQNHDV0 ( QN, CK, D, E, VDD, VSS); 
input CK, D, E;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  not      I1 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_E,dE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            negedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            posedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK, posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDQNHDV2 ( QN, CK, D, E, VDD, VSS); 
input CK, D, E;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  not      I1 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_E,dE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            negedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            posedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK, posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDQNHDV4 ( QN, CK, D, E, VDD, VSS); 
input CK, D, E;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  not      I1 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_E,dE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            negedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            posedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK, posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDQNHDV8 ( QN, CK, D, E, VDD, VSS); 
input CK, D, E;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  not      I1 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    buf SMC_I6(ENABLE_E,dE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            negedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E === 1'b1), 
            posedge D &&& (ENABLE_E === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
        $setuphold(posedge CK, posedge E, 1.0, 1.0, NOTIFIER, , , dCK, dE); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDRNQHDV0 (D, E, RDN, CK, Q, VDD, VSS); 
  input D, E, RDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_E;
  buf    XX0 (xRN, dRDN );
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  buf     B1 (Q_temp, n0 );
  assign ENABLE_D_AND_E = ( D & E )?1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(ENABLE_E_AND_RDN,dE,dRDN);

    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1), posedge RDN &&& (ENABLE_D_AND_E === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDRNQHDV2 (D, E, RDN, CK, Q, VDD, VSS); 
  input D, E, RDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_E;
  buf    XX0 (xRN, dRDN );
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  buf     B1 (Q_temp, n0 );
  assign ENABLE_D_AND_E = ( D & E )?1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(ENABLE_E_AND_RDN,dE,dRDN);

    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1), posedge RDN &&& (ENABLE_D_AND_E === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDRNQHDV4 (D, E, RDN, CK, Q, VDD, VSS); 
  input D, E, RDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_E;
  buf    XX0 (xRN, dRDN );
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  buf     B1 (Q_temp, n0 );
  assign ENABLE_D_AND_E = ( D & E )?1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(ENABLE_E_AND_RDN,dE,dRDN);

    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1), posedge RDN &&& (ENABLE_D_AND_E === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDRNQHDV8 (D, E, RDN, CK, Q, VDD, VSS); 
  input D, E, RDN, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_E;
  buf    XX0 (xRN, dRDN );
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  buf     B1 (Q_temp, n0 );
  assign ENABLE_D_AND_E = ( D & E )?1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(ENABLE_E_AND_RDN,dE,dRDN);

    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1), posedge RDN &&& (ENABLE_D_AND_E === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDRNQNHDV0 (D, E, RDN, CK, QN, VDD, VSS); 
  input D, E, RDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_E;
  buf     XX0 (xRN, dRDN );
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  not      I1 (QN_temp, n0 );
  assign ENABLE_D_AND_E = ( D & E )?1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_E_AND_RDN,dE,dRDN);

    buf SMC_I7(ENABLE_RDN,dRDN);


  specify


	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1), posedge RDN &&& (ENABLE_D_AND_E === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDRNQNHDV2 (D, E, RDN, CK, QN, VDD, VSS); 
  input D, E, RDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_E;
  buf     XX0 (xRN, dRDN );
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  not      I1 (QN_temp, n0 );
  assign ENABLE_D_AND_E = ( D & E )?1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_E_AND_RDN,dE,dRDN);

    buf SMC_I7(ENABLE_RDN,dRDN);


  specify


	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1), posedge RDN &&& (ENABLE_D_AND_E === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDRNQNHDV4 (D, E, RDN, CK, QN, VDD, VSS); 
  input D, E, RDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_E;
  buf     XX0 (xRN, dRDN );
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  not      I1 (QN_temp, n0 );
  assign ENABLE_D_AND_E = ( D & E )?1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_E_AND_RDN,dE,dRDN);

    buf SMC_I7(ENABLE_RDN,dRDN);


  specify


	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1), posedge RDN &&& (ENABLE_D_AND_E === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module EDRNQNHDV8 (D, E, RDN, CK, QN, VDD, VSS); 
  input D, E, RDN, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_E;
  buf     XX0 (xRN, dRDN );
  udp_edff_PWR I0 (n0, dD, dCK, xRN, xSN, dE, VDD, VSS, NOTIFIER ); 
  not      I1 (QN_temp, n0 );
  assign ENABLE_D_AND_E = ( D & E )?1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_E_AND_RDN,dE,dRDN);

    buf SMC_I7(ENABLE_RDN,dRDN);


  specify


	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge E &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E === 1'b1), posedge RDN &&& (ENABLE_D_AND_E === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHHDV0 ( Q, QN, D, E, VDD, VSS); 
input D, E;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  not I3(clk, dE );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc D --> Q 
	 (D => Q) = (1.0,1.0); 
 
	// arc E --> Q 
	(posedge E => (Q : D))  = (1.0,1.0); 
 
	// arc D --> QN 
	 (D => QN) = (1.0,1.0); 
 
	// arc E --> QN 
	(posedge E => (QN : D))  = (1.0,1.0); 
 
        $setuphold(negedge E, negedge D, 1.0, 1.0, NOTIFIER, , , dE, dD); 
 
        $setuphold(negedge E, posedge D, 1.0, 1.0, NOTIFIER, , , dE, dD); 
 
 
 
        $width(posedge E,1.0,0,NOTIFIER); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHHDV2 ( Q, QN, D, E, VDD, VSS); 
input D, E;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  not I3(clk, dE );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc D --> Q 
	 (D => Q) = (1.0,1.0); 
 
	// arc E --> Q 
	(posedge E => (Q : D))  = (1.0,1.0); 
 
	// arc D --> QN 
	 (D => QN) = (1.0,1.0); 
 
	// arc E --> QN 
	(posedge E => (QN : D))  = (1.0,1.0); 
 
        $setuphold(negedge E, negedge D, 1.0, 1.0, NOTIFIER, , , dE, dD); 
 
        $setuphold(negedge E, posedge D, 1.0, 1.0, NOTIFIER, , , dE, dD); 
 
 
 
        $width(posedge E,1.0,0,NOTIFIER); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHHDV4 ( Q, QN, D, E, VDD, VSS); 
input D, E;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  not I3(clk, dE );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc D --> Q 
	 (D => Q) = (1.0,1.0); 
 
	// arc E --> Q 
	(posedge E => (Q : D))  = (1.0,1.0); 
 
	// arc D --> QN 
	 (D => QN) = (1.0,1.0); 
 
	// arc E --> QN 
	(posedge E => (QN : D))  = (1.0,1.0); 
 
        $setuphold(negedge E, negedge D, 1.0, 1.0, NOTIFIER, , , dE, dD); 
 
        $setuphold(negedge E, posedge D, 1.0, 1.0, NOTIFIER, , , dE, dD); 
 
 
 
        $width(posedge E,1.0,0,NOTIFIER); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHRNHDV0 (D, RDN, E, Q, QN, VDD, VSS); 
  input D, RDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
not      I3(clk, dE );
buf      XX0 (xRN, dRDN );
udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
buf      I1 (Q_temp, n0 );
not      I2 (QN_temp, n0 );
assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dE, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHRNHDV2 (D, RDN, E, Q, QN, VDD, VSS); 
  input D, RDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
not      I3(clk, dE );
buf      XX0 (xRN, dRDN );
udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
buf      I1 (Q_temp, n0 );
not      I2 (QN_temp, n0 );
assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dE, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHRNHDV4 (D, RDN, E, Q, QN, VDD, VSS); 
  input D, RDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
not      I3(clk, dE );
buf      XX0 (xRN, dRDN );
udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
buf      I1 (Q_temp, n0 );
not      I2 (QN_temp, n0 );
assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_RDN,dRDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dE, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHRSNHDV0 (D, RDN, SDN, E, Q, QN, VDD, VSS); 
  input D, RDN, SDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf       XX0 (xSN, dSDN );
  buf       XX1 (xRN, dRDN );
  not I3(clk, dE );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);
    
    not SMC_I9(ENABLE_NOT_E,dE);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dSDN);


        $setuphold(posedge RDN &&& (ENABLE_NOT_E === 1'b1),
            posedge SDN &&& (ENABLE_NOT_E === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHRSNHDV2 (D, RDN, SDN, E, Q, QN, VDD, VSS); 
  input D, RDN, SDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf       XX0 (xSN, dSDN );
  buf       XX1 (xRN, dRDN );
  not I3(clk, dE );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);
    
    not SMC_I9(ENABLE_NOT_E,dE);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dSDN);


        $setuphold(posedge RDN &&& (ENABLE_NOT_E === 1'b1),
            posedge SDN &&& (ENABLE_NOT_E === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHRSNHDV4 (D, RDN, SDN, E, Q, QN, VDD, VSS); 
  input D, RDN, SDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf       XX0 (xSN, dSDN );
  buf       XX1 (xRN, dRDN );
  not I3(clk, dE );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I7(ENABLE_SDN,dSDN);

    buf SMC_I8(ENABLE_RDN,dRDN);
    
    not SMC_I9(ENABLE_NOT_E,dE);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dSDN);


        $setuphold(posedge RDN &&& (ENABLE_NOT_E === 1'b1),
            posedge SDN &&& (ENABLE_NOT_E === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHSNHDV0 (D, SDN, E, Q, QN, VDD, VSS); 
  input D, SDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  not      I3 (clk, dE );
  buf      XX0 (xSN, dSDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dE, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHSNHDV2 (D, SDN, E, Q, QN, VDD, VSS); 
  input D, SDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  not      I3 (clk, dE );
  buf      XX0 (xSN, dSDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dE, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LAHSNHDV4 (D, SDN, E, Q, QN, VDD, VSS); 
  input D, SDN, E;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  not      I3 (clk, dE );
  buf      XX0 (xSN, dSDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc E --> Q
	(posedge E => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc E --> QN
	(posedge E => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && E===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && E===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && E===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(negedge E &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);

        $setuphold(negedge E &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dE, dD);



        $width(posedge E,1.0,0,NOTIFIER);

        $setuphold(negedge E &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dE, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALHDV0 ( Q, QN, D, EN, VDD, VSS); 
input D, EN;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf      I3 (clk, dEN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc D --> Q 
	 (D => Q) = (1.0,1.0); 
 
	// arc EN --> Q 
	(negedge EN => (Q : D))  = (1.0,1.0); 
 
	// arc D --> QN 
	 (D => QN) = (1.0,1.0); 
 
	// arc EN --> QN 
	(negedge EN => (QN : D))  = (1.0,1.0); 
 
        $setuphold(posedge EN, negedge D, 1.0, 1.0, NOTIFIER, , , dEN, dD); 
 
        $setuphold(posedge EN, posedge D, 1.0, 1.0, NOTIFIER, , , dEN, dD); 
 
 
 
        $width(negedge EN,1.0,0,NOTIFIER); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALHDV2 ( Q, QN, D, EN, VDD, VSS); 
input D, EN;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf      I3 (clk, dEN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc D --> Q 
	 (D => Q) = (1.0,1.0); 
 
	// arc EN --> Q 
	(negedge EN => (Q : D))  = (1.0,1.0); 
 
	// arc D --> QN 
	 (D => QN) = (1.0,1.0); 
 
	// arc EN --> QN 
	(negedge EN => (QN : D))  = (1.0,1.0); 
 
        $setuphold(posedge EN, negedge D, 1.0, 1.0, NOTIFIER, , , dEN, dD); 
 
        $setuphold(posedge EN, posedge D, 1.0, 1.0, NOTIFIER, , , dEN, dD); 
 
 
 
        $width(negedge EN,1.0,0,NOTIFIER); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALHDV4 ( Q, QN, D, EN, VDD, VSS); 
input D, EN;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf      I3 (clk, dEN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc D --> Q 
	 (D => Q) = (1.0,1.0); 
 
	// arc EN --> Q 
	(negedge EN => (Q : D))  = (1.0,1.0); 
 
	// arc D --> QN 
	 (D => QN) = (1.0,1.0); 
 
	// arc EN --> QN 
	(negedge EN => (QN : D))  = (1.0,1.0); 
 
        $setuphold(posedge EN, negedge D, 1.0, 1.0, NOTIFIER, , , dEN, dD); 
 
        $setuphold(posedge EN, posedge D, 1.0, 1.0, NOTIFIER, , , dEN, dD); 
 
 
 
        $width(negedge EN,1.0,0,NOTIFIER); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALRNHDV0 (D, RDN, EN, Q, QN, VDD, VSS); 
  input D, RDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf      I3 (clk, dEN );
  buf       XX0 (xRN, dRDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_RDN,dRDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dEN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALRNHDV2 (D, RDN, EN, Q, QN, VDD, VSS); 
  input D, RDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf      I3 (clk, dEN );
  buf       XX0 (xRN, dRDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_RDN,dRDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dEN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALRNHDV4 (D, RDN, EN, Q, QN, VDD, VSS); 
  input D, RDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf      I3 (clk, dEN );
  buf       XX0 (xRN, dRDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_RDN,dRDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dEN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALRSNHDV0 (D, RDN, SDN, EN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf      I3 (clk, dEN );
  buf      XX0 (xSN, dSDN );
  buf      XX1 (xRN, dRDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I8(ENABLE_SDN,dSDN);

    buf SMC_I9(ENABLE_RDN,dRDN);

    buf SMC_I10(ENABLE_EN,dEN);

  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dSDN);


        $setuphold(posedge RDN &&& (ENABLE_EN === 1'b1),
            posedge SDN &&& (ENABLE_EN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALRSNHDV2 (D, RDN, SDN, EN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf      I3 (clk, dEN );
  buf      XX0 (xSN, dSDN );
  buf      XX1 (xRN, dRDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I8(ENABLE_SDN,dSDN);

    buf SMC_I9(ENABLE_RDN,dRDN);

    buf SMC_I10(ENABLE_EN,dEN);

  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dSDN);


        $setuphold(posedge RDN &&& (ENABLE_EN === 1'b1),
            posedge SDN &&& (ENABLE_EN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALRSNHDV4 (D, RDN, SDN, EN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf      I3 (clk, dEN );
  buf      XX0 (xSN, dSDN );
  buf      XX1 (xRN, dRDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I8(ENABLE_SDN,dSDN);

    buf SMC_I9(ENABLE_RDN,dRDN);

    buf SMC_I10(ENABLE_EN,dEN);

  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dSDN);


        $setuphold(posedge RDN &&& (ENABLE_EN === 1'b1),
            posedge SDN &&& (ENABLE_EN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALSNHDV0 (D, SDN, EN, Q, QN, VDD, VSS); 
  input D, SDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf      I3 (clk, dEN );
  buf      XX0 (xSN, dSDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_SDN,dSDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dEN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALSNHDV2 (D, SDN, EN, Q, QN, VDD, VSS); 
  input D, SDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf      I3 (clk, dEN );
  buf      XX0 (xSN, dSDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_SDN,dSDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dEN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module LALSNHDV4 (D, SDN, EN, Q, QN, VDD, VSS); 
  input D, SDN, EN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf      I3 (clk, dEN );
  buf      XX0 (xSN, dSDN );
  udp_tlat_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf      I1 (Q_temp, n0 );
  not      I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_SDN,dSDN);


  specify


	// arc D --> Q
	 (D => Q) = (1.0,1.0);

	// arc EN --> Q
	(negedge EN => (Q : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc D --> QN
	 (D => QN) = (1.0,1.0);

	// arc EN --> QN
	(negedge EN => (QN : D))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b0 && EN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(D===1'b1 && EN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $setuphold(posedge EN &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);

        $setuphold(posedge EN &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dEN, dD);



        $width(negedge EN,1.0,0,NOTIFIER);

        $setuphold(posedge EN &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dEN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2HDV0 ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2HDV1 ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2HDV2 ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2HDV4 ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2HDVL ( Z, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux2_PWR (Z_temp, I0, I1, S ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 

        if(I1===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

 	ifnone
	(I0 => Z) = (1.0,1.0);	
  
	if(I0===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

 	ifnone
	(I1 => Z) = (1.0,1.0);	
 
	// arc posedge S --> (Z:S) 
	 (posedge S => (Z:S)) = (1.0,1.0); 
 
	// arc negedge S --> (Z:S) 
	 (negedge S => (Z:S)) = (1.0,1.0);
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2NHDV0 ( ZN, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  udp_mux2_PWR I00(z, I0, I1, S ,VDD, VSS); 
  not      I01(ZN_temp, z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 	
	ifnone
	(I0 => ZN) = (1.0,1.0);	
 
	if(I0===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	(I1 => ZN) = (1.0,1.0);	
 
	// arc posedge S --> (ZN:S) 
	 (posedge S => (ZN:S)) = (1.0,1.0); 
 
	// arc negedge S --> (ZN:S) 
	 (negedge S => (ZN:S)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2NHDV1 ( ZN, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  udp_mux2_PWR I00(z, I0, I1, S ,VDD, VSS); 
  not      I01(ZN_temp, z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 	
	ifnone
	(I0 => ZN) = (1.0,1.0);	
 
	if(I0===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	(I1 => ZN) = (1.0,1.0);	
 
	// arc posedge S --> (ZN:S) 
	 (posedge S => (ZN:S)) = (1.0,1.0); 
 
	// arc negedge S --> (ZN:S) 
	 (negedge S => (ZN:S)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2NHDV2 ( ZN, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  udp_mux2_PWR I00(z, I0, I1, S ,VDD, VSS); 
  not      I01(ZN_temp, z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 	
	ifnone
	(I0 => ZN) = (1.0,1.0);	
 
	if(I0===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	(I1 => ZN) = (1.0,1.0);	
 
	// arc posedge S --> (ZN:S) 
	 (posedge S => (ZN:S)) = (1.0,1.0); 
 
	// arc negedge S --> (ZN:S) 
	 (negedge S => (ZN:S)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2NHDV4 ( ZN, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  udp_mux2_PWR I00(z, I0, I1, S ,VDD, VSS); 
  not      I01(ZN_temp, z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 	
	ifnone
	(I0 => ZN) = (1.0,1.0);	
 
	if(I0===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	(I1 => ZN) = (1.0,1.0);	
 
	// arc posedge S --> (ZN:S) 
	 (posedge S => (ZN:S)) = (1.0,1.0); 
 
	// arc negedge S --> (ZN:S) 
	 (negedge S => (ZN:S)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX2NHDVL ( ZN, I0, I1, S, VDD, VSS); 
input I0, I1, S;
inout VDD, VSS;
output ZN;
wire ZN_temp;

  udp_mux2_PWR I00(z, I0, I1, S ,VDD, VSS); 
  not      I01(ZN_temp, z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 	
	ifnone
	(I0 => ZN) = (1.0,1.0);	
 
	if(I0===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	(I1 => ZN) = (1.0,1.0);	
 
	// arc posedge S --> (ZN:S) 
	 (posedge S => (ZN:S)) = (1.0,1.0); 
 
	// arc negedge S --> (ZN:S) 
	 (negedge S => (ZN:S)) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3HDV0 ( Z, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux4_PWR u0 (Z_temp, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

	ifnone
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

	ifnone
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 

	ifnone
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3HDV1 ( Z, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux4_PWR u0 (Z_temp, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

	ifnone
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

	ifnone
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 

	ifnone
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3HDV2 ( Z, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux4_PWR u0 (Z_temp, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

	ifnone
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

	ifnone
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 

	ifnone
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3HDV4 ( Z, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux4_PWR u0 (Z_temp, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

	ifnone
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

	ifnone
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 

	ifnone
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3HDVL ( Z, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output Z;
wire Z_temp;

  udp_mux4_PWR u0 (Z_temp, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
  assign Z = ((VDD === 1'b1) && (VSS === 1'b0)) ? Z_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 

	ifnone
	// arc I0 --> Z 
	 (I0 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 

	ifnone
	// arc I1 --> Z 
	 (I1 => Z) = (1.0,1.0); 




 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 

	ifnone
	// arc I2 --> Z 
	 (I2 => Z) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (Z:S0) 
	 (posedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (Z:S0) 
	 (negedge S0 => (Z:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> Z 
	 (S1 => Z) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3NHDV0 ( ZN, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   udp_mux4_PWR u0 (Z, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
   not u1(ZN_temp, Z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 

	ifnone 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 


 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 



 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 

	ifnone
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3NHDV1 ( ZN, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   udp_mux4_PWR u0 (Z, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
   not u1(ZN_temp, Z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 

	ifnone 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 


 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 



 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 

	ifnone
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3NHDV2 ( ZN, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   udp_mux4_PWR u0 (Z, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
   not u1(ZN_temp, Z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 

	ifnone 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 


 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 



 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 

	ifnone
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3NHDV4 ( ZN, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   udp_mux4_PWR u0 (Z, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
   not u1(ZN_temp, Z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 

	ifnone 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 


 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 



 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 

	ifnone
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module MUX3NHDVL ( ZN, I0, I1, I2, S0, S1, VDD, VSS); 
input I0, I1, I2, S0, S1;
inout VDD, VSS;
output ZN;
wire ZN_temp;

   udp_mux4_PWR u0 (Z, I0, I1, I2, I2, S0, S1 ,VDD, VSS); 
   not u1(ZN_temp, Z );
  assign ZN = ((VDD === 1'b1) && (VSS === 1'b0)) ? ZN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	if(I1===1'b0 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b0 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b0) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 
 
	if(I1===1'b1 && I2===1'b1) 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 

	ifnone 
	// arc I0 --> ZN 
	 (I0 => ZN) = (1.0,1.0); 


 
	if(I0===1'b0 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b0) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I2===1'b1) 
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 

	ifnone
	// arc I1 --> ZN 
	 (I1 => ZN) = (1.0,1.0); 



 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 

	ifnone
	// arc I2 --> ZN 
	 (I2 => ZN) = (1.0,1.0); 




 
	if(I2===1'b0) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b0) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc posedge S0 --> (ZN:S0) 
	 (posedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I2===1'b1) 
	// arc negedge S0 --> (ZN:S0) 
	 (negedge S0 => (ZN:S0)) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b0 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b0 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b0) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
	if(I0===1'b1 && I1===1'b1 && S0===1'b1) 
	// arc S1 --> ZN 
	 (S1 => ZN) = (1.0,1.0); 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDHDV0 ( Q, QN, CKN, D, VDD, VSS); 
input CKN, D;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CKN --> Q 
	(negedge CKN => (Q : D))  = (1.0,1.0); 
 
	// arc CKN --> QN 
	(negedge CKN => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CKN,1.0,0,NOTIFIER); 
 
        $width(posedge CKN,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CKN, negedge D, 1.0, 1.0, NOTIFIER, , , dCKN, dD); 
 
        $setuphold(negedge CKN, posedge D, 1.0, 1.0, NOTIFIER, , , dCKN, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDHDV2 ( Q, QN, CKN, D, VDD, VSS); 
input CKN, D;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CKN --> Q 
	(negedge CKN => (Q : D))  = (1.0,1.0); 
 
	// arc CKN --> QN 
	(negedge CKN => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CKN,1.0,0,NOTIFIER); 
 
        $width(posedge CKN,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CKN, negedge D, 1.0, 1.0, NOTIFIER, , , dCKN, dD); 
 
        $setuphold(negedge CKN, posedge D, 1.0, 1.0, NOTIFIER, , , dCKN, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDHDV4 ( Q, QN, CKN, D, VDD, VSS); 
input CKN, D;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN,xRN; 
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
 
  specify 
 
 
	// arc CKN --> Q 
	(negedge CKN => (Q : D))  = (1.0,1.0); 
 
	// arc CKN --> QN 
	(negedge CKN => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CKN,1.0,0,NOTIFIER); 
 
        $width(posedge CKN,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CKN, negedge D, 1.0, 1.0, NOTIFIER, , , dCKN, dD); 
 
        $setuphold(negedge CKN, posedge D, 1.0, 1.0, NOTIFIER, , , dCKN, dD); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDRNHDV0 (D, RDN, CKN, Q, QN, VDD, VSS); 
  input D, RDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_RDN,dRDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDRNHDV2 (D, RDN, CKN, Q, QN, VDD, VSS); 
  input D, RDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_RDN,dRDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDRNHDV4 (D, RDN, CKN, Q, QN, VDD, VSS); 
  input D, RDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D;
  buf   XX0 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_D= (D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(ENABLE_RDN,dRDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            negedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            posedge D &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D === 1'b1), posedge RDN &&& (ENABLE_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDRSNHDV0 (D, RDN, SDN, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I8(ENABLE_SDN,dSDN);

    buf SMC_I9(ENABLE_RDN,dRDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDRSNHDV2 (D, RDN, SDN, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I8(ENABLE_SDN,dSDN);

    buf SMC_I9(ENABLE_RDN,dRDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDRSNHDV4 (D, RDN, SDN, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN;
wire ENABLE_NOT_D_AND_RDN;
  buf   XX0 (xSN, dSDN );
  buf   XX1 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN = ( D & SDN )? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN = ( !D & RDN ) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    and SMC_I7(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    buf SMC_I8(ENABLE_SDN,dSDN);

    buf SMC_I9(ENABLE_RDN,dRDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_SDN === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_RDN === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDSNHDV0 (D, SDN, CKN, Q, QN, VDD, VSS); 
  input D, SDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDSNHDV2 (D, SDN, CKN, Q, QN, VDD, VSS); 
  input D, SDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module NDSNHDV4 (D, SDN, CKN, Q, QN, VDD, VSS); 
  input D, SDN, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D;
  buf   XX0 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, dD, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  not     I2 (QN_temp, n0 );
  assign ENABLE_NOT_D= (!D) ? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(ENABLE_SDN,dSDN);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            negedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            posedge D &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_NOT_D === 1'b1), posedge SDN &&& (ENABLE_NOT_D === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);


  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDGRNQHDV0 ( Q, CK, D, RN, SE, SI, VDD, VSS); 
input CK, D, RN, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN; 
  buf   XX0 (xRN, dRN );
  udp_sedfft_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER ); 
  buf        I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I7(ENABLE_NOT_SE,dSE); 
 
 
    buf SMC_I9(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDGRNQHDV2 ( Q, CK, D, RN, SE, SI, VDD, VSS); 
input CK, D, RN, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN; 
  buf   XX0 (xRN, dRN );
  udp_sedfft_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER ); 
  buf        I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I7(ENABLE_NOT_SE,dSE); 
 
 
    buf SMC_I9(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDGRNQHDV4 ( Q, CK, D, RN, SE, SI, VDD, VSS); 
input CK, D, RN, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN; 
  buf   XX0 (xRN, dRN );
  udp_sedfft_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER ); 
  buf        I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I7(ENABLE_NOT_SE,dSE); 
 
 
    buf SMC_I9(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDGRNQHDV8 ( Q, CK, D, RN, SE, SI, VDD, VSS); 
input CK, D, RN, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xSN; 
  buf   XX0 (xRN, dRN );
  udp_sedfft_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER ); 
  buf        I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I7(ENABLE_NOT_SE,dSE); 
 
 
    buf SMC_I9(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDGRNQNHDV0 ( QN, CK, D, RN, SE, SI, VDD, VSS); 
input CK, D, RN, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN; 
  buf   XX0 (xRN, dRN );
  udp_sedfft_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER ); 
  not        I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I10(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I11(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDGRNQNHDV2 ( QN, CK, D, RN, SE, SI, VDD, VSS); 
input CK, D, RN, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN; 
  buf   XX0 (xRN, dRN );
  udp_sedfft_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER ); 
  not        I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I10(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I11(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDGRNQNHDV4 ( QN, CK, D, RN, SE, SI, VDD, VSS); 
input CK, D, RN, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN; 
  buf   XX0 (xRN, dRN );
  udp_sedfft_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER ); 
  not        I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I10(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I11(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDGRNQNHDV8 ( QN, CK, D, RN, SE, SI, VDD, VSS); 
input CK, D, RN, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xSN; 
  buf   XX0 (xRN, dRN );
  udp_sedfft_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, 1'b1, VDD, VSS, NOTIFIER ); 
  not        I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I10(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I11(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge RN &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dRN); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDQHDV0 ( Q, CK, D, SE, SI, VDD, VSS); 
input CK, D, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I4(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I5(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDQHDV2 ( Q, CK, D, SE, SI, VDD, VSS); 
input CK, D, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I4(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I5(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDQHDV4 ( Q, CK, D, SE, SI, VDD, VSS); 
input CK, D, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I4(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I5(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDQHDV8 ( Q, CK, D, SE, SI, VDD, VSS); 
input CK, D, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I4(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I5(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDQNHDV0 ( QN, CK, D, SE, SI, VDD, VSS); 
input CK, D, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I6(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I7(ENABLE_SE,dSE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDQNHDV2 ( QN, CK, D, SE, SI, VDD, VSS); 
input CK, D, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I6(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I7(ENABLE_SE,dSE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDQNHDV4 ( QN, CK, D, SE, SI, VDD, VSS); 
input CK, D, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I6(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I7(ENABLE_SE,dSE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDQNHDV8 ( QN, CK, D, SE, SI, VDD, VSS); 
input CK, D, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I6(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I7(ENABLE_SE,dSE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRNQHDV0 (D, RDN, SE, SI, CK, Q, VDD, VSS); 
  input D, RDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I6(ENABLE_RDN,dRDN);

    and SMC_I7(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRNQHDV2 (D, RDN, SE, SI, CK, Q, VDD, VSS); 
  input D, RDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I6(ENABLE_RDN,dRDN);

    and SMC_I7(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRNQHDV4 (D, RDN, SE, SI, CK, Q, VDD, VSS); 
  input D, RDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I6(ENABLE_RDN,dRDN);

    and SMC_I7(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRNQHDV8 (D, RDN, SE, SI, CK, Q, VDD, VSS); 
  input D, RDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I6(ENABLE_RDN,dRDN);

    and SMC_I7(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRNQNHDV0 (D, RDN, SE, SI, CK, QN, VDD, VSS); 
  input D, RDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional
				// none
  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I8(ENABLE_RDN,dRDN);

    and SMC_I9(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRNQNHDV2 (D, RDN, SE, SI, CK, QN, VDD, VSS); 
  input D, RDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional
				// none
  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I8(ENABLE_RDN,dRDN);

    and SMC_I9(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRNQNHDV4 (D, RDN, SE, SI, CK, QN, VDD, VSS); 
  input D, RDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional
				// none
  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I8(ENABLE_RDN,dRDN);

    and SMC_I9(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRNQNHDV8 (D, RDN, SE, SI, CK, QN, VDD, VSS); 
  input D, RDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional
				// none
  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I8(ENABLE_RDN,dRDN);

    and SMC_I9(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRQHDV0 (D, RD, SE, SI, CK, Q, VDD, VSS); 
  input D, RD, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_NOT_RD_AND_NOT_SE,xRN, SE_bar);

    not SMC_I6(ENABLE_NOT_RD,dRD);

    and SMC_I7(ENABLE_NOT_RD_AND_SE,xRN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), negedge RD &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRQHDV2 (D, RD, SE, SI, CK, Q, VDD, VSS); 
  input D, RD, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_NOT_RD_AND_NOT_SE,xRN, SE_bar);

    not SMC_I6(ENABLE_NOT_RD,dRD);

    and SMC_I7(ENABLE_NOT_RD_AND_SE,xRN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), negedge RD &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRQHDV4 (D, RD, SE, SI, CK, Q, VDD, VSS); 
  input D, RD, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_NOT_RD_AND_NOT_SE,xRN, SE_bar);

    not SMC_I6(ENABLE_NOT_RD,dRD);

    and SMC_I7(ENABLE_NOT_RD_AND_SE,xRN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), negedge RD &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRQHDV8 (D, RD, SE, SI, CK, Q, VDD, VSS); 
  input D, RD, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_NOT_RD_AND_NOT_SE,xRN, SE_bar);

    not SMC_I6(ENABLE_NOT_RD,dRD);

    and SMC_I7(ENABLE_NOT_RD_AND_SE,xRN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> Q
	(posedge RD => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), negedge RD &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRQNHDV0 (D, RD, SE, SI, CK, QN, VDD, VSS); 
  input D, RD, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional
				// none
  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_NOT_RD_AND_NOT_SE,xRN, SE_bar);

    not SMC_I8(ENABLE_NOT_RD,dRD);

    and SMC_I9(ENABLE_NOT_RD_AND_SE,xRN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), negedge RD &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRQNHDV2 (D, RD, SE, SI, CK, QN, VDD, VSS); 
  input D, RD, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional
				// none
  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_NOT_RD_AND_NOT_SE,xRN, SE_bar);

    not SMC_I8(ENABLE_NOT_RD,dRD);

    and SMC_I9(ENABLE_NOT_RD_AND_SE,xRN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), negedge RD &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRQNHDV4 (D, RD, SE, SI, CK, QN, VDD, VSS); 
  input D, RD, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional
				// none
  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_NOT_RD_AND_NOT_SE,xRN, SE_bar);

    not SMC_I8(ENABLE_NOT_RD,dRD);

    and SMC_I9(ENABLE_NOT_RD_AND_SE,xRN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), negedge RD &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRQNHDV8 (D, RD, SE, SI, CK, QN, VDD, VSS); 
  input D, RD, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  not   XX0 (xRN, dRD );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional
				// none
  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_NOT_RD_AND_NOT_SE,xRN, SE_bar);

    not SMC_I8(ENABLE_NOT_RD,dRD);

    and SMC_I9(ENABLE_NOT_RD_AND_SE,xRN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RD --> QN
	(posedge RD => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_NOT_RD_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), negedge RD &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRD);


        $width(posedge RD,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            negedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD === 1'b1),
            posedge SE &&& (ENABLE_NOT_RD === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_NOT_RD_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_NOT_RD_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRSNQHDV0 (D, RDN, SDN, SE, SI, CK, Q, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);

    and SMC_I8(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    buf SMC_I10(ENABLE_RDN,dRDN);

    and SMC_I11(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I12(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	
        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRSNQHDV2 (D, RDN, SDN, SE, SI, CK, Q, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);

    and SMC_I8(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    buf SMC_I10(ENABLE_RDN,dRDN);

    and SMC_I11(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I12(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	
        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRSNQHDV4 (D, RDN, SDN, SE, SI, CK, Q, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);

    and SMC_I8(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    buf SMC_I10(ENABLE_RDN,dRDN);

    and SMC_I11(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I12(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	
        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRSNQHDV8 (D, RDN, SDN, SE, SI, CK, Q, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);

    and SMC_I8(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    buf SMC_I10(ENABLE_RDN,dRDN);

    and SMC_I11(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I12(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	
        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRSNQNHDV0 (D, RDN, SDN, SE, SI, CK, QN, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CK;
inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);

    and SMC_I8(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    buf SMC_I10(ENABLE_RDN,dRDN);

    and SMC_I11(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I12(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRSNQNHDV2 (D, RDN, SDN, SE, SI, CK, QN, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CK;
inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);

    and SMC_I8(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    buf SMC_I10(ENABLE_RDN,dRDN);

    and SMC_I11(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I12(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRSNQNHDV4 (D, RDN, SDN, SE, SI, CK, QN, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CK;
inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);

    and SMC_I8(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    buf SMC_I10(ENABLE_RDN,dRDN);

    and SMC_I11(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I12(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDRSNQNHDV8 (D, RDN, SDN, SE, SI, CK, QN, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CK;
inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);

    and SMC_I8(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    buf SMC_I10(ENABLE_RDN,dRDN);

    and SMC_I11(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I12(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDSNQHDV0 (D, SDN, SE, SI, CK, Q, VDD, VSS); 
  input D, SDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);

    and SMC_I7(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I8(ENABLE_SDN,dSDN);

    and SMC_I9(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);


        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDSNQHDV2 (D, SDN, SE, SI, CK, Q, VDD, VSS); 
  input D, SDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);

    and SMC_I7(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I8(ENABLE_SDN,dSDN);

    and SMC_I9(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);


        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDSNQHDV4 (D, SDN, SE, SI, CK, Q, VDD, VSS); 
  input D, SDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);

    and SMC_I7(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I8(ENABLE_SDN,dSDN);

    and SMC_I9(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);


        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDSNQHDV8 (D, SDN, SE, SI, CK, Q, VDD, VSS); 
  input D, SDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);

    and SMC_I7(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I8(ENABLE_SDN,dSDN);

    and SMC_I9(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);


        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDSNQNHDV0 (D, SDN, SE, SI, CK, QN, VDD, VSS); 
  input D, SDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);

    and SMC_I7(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I8(ENABLE_SDN,dSDN);

    and SMC_I9(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDSNQNHDV2 (D, SDN, SE, SI, CK, QN, VDD, VSS); 
  input D, SDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);

    and SMC_I7(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I8(ENABLE_SDN,dSDN);

    and SMC_I9(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDSNQNHDV4 (D, SDN, SE, SI, CK, QN, VDD, VSS); 
  input D, SDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);

    and SMC_I7(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I8(ENABLE_SDN,dSDN);

    and SMC_I9(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDSNQNHDV8 (D, SDN, SE, SI, CK, QN, VDD, VSS); 
  input D, SDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  not     I3 (QN_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);

    and SMC_I7(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I8(ENABLE_SDN,dSDN);

    and SMC_I9(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDXHDV0 ( Q, QN, CK, DA, DB, SA, SE, SI, VDD, VSS); 
input CK, DA, DB, SA, SE, SI;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n2, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n2, n1, dSI, dSE ,VDD, VSS); 
  udp_mux_PWR I2 (n1, dDB, dDA, dSA ,VDD, VSS); 
  buf     I3 (Q_temp, n0 );
  not     I4 (QN_temp, n0 );
  not     I5 (SE_bar, dSE );
  not     I6 (SA_bar, dSA );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    and SMC_I11(ENABLE_SA_AND_NOT_SE,dSA, SE_bar); 
 
    and SMC_I12(ENABLE_NOT_SA_AND_NOT_SE, SA_bar, SE_bar); 
 
    not SMC_I13(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I14(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : DA))  = (1.0,1.0); 
 
	// arc CK --> QN 
	(posedge CK => (QN : DA))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 
            negedge DA &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
        $setuphold(posedge CK &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 
            posedge DA &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 
            negedge DB &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 
            posedge DB &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge SA &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSA); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge SA &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSA); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDXHDV2 ( Q, QN, CK, DA, DB, SA, SE, SI, VDD, VSS); 
input CK, DA, DB, SA, SE, SI;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n2, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n2, n1, dSI, dSE ,VDD, VSS); 
  udp_mux_PWR I2 (n1, dDB, dDA, dSA ,VDD, VSS); 
  buf     I3 (Q_temp, n0 );
  not     I4 (QN_temp, n0 );
  not     I5 (SE_bar, dSE );
  not     I6 (SA_bar, dSA );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    and SMC_I11(ENABLE_SA_AND_NOT_SE,dSA, SE_bar); 
 
    and SMC_I12(ENABLE_NOT_SA_AND_NOT_SE, SA_bar, SE_bar); 
 
    not SMC_I13(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I14(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : DA))  = (1.0,1.0); 
 
	// arc CK --> QN 
	(posedge CK => (QN : DA))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 
            negedge DA &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
        $setuphold(posedge CK &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 
            posedge DA &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 
            negedge DB &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 
            posedge DB &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge SA &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSA); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge SA &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSA); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SDXHDV4 ( Q, QN, CK, DA, DB, SA, SE, SI, VDD, VSS); 
input CK, DA, DB, SA, SE, SI;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  buf     IC (clk, dCK );
  udp_dff_PWR I0 (n0, n2, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n2, n1, dSI, dSE ,VDD, VSS); 
  udp_mux_PWR I2 (n1, dDB, dDA, dSA ,VDD, VSS); 
  buf     I3 (Q_temp, n0 );
  not     I4 (QN_temp, n0 );
  not     I5 (SE_bar, dSE );
  not     I6 (SA_bar, dSA );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    and SMC_I11(ENABLE_SA_AND_NOT_SE,dSA, SE_bar); 
 
    and SMC_I12(ENABLE_NOT_SA_AND_NOT_SE, SA_bar, SE_bar); 
 
    not SMC_I13(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I14(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : DA))  = (1.0,1.0); 
 
	// arc CK --> QN 
	(posedge CK => (QN : DA))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 
            negedge DA &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
        $setuphold(posedge CK &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 
            posedge DA &&& (ENABLE_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDA); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 
            negedge DB &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 
            posedge DB &&& (ENABLE_NOT_SA_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dDB); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge SA &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSA); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge SA &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSA); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDQHDV0 ( Q, CK, D, E, SE, SI, VDD, VSS); 
input CK, D, E, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_sedff_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I4(SE_bar,dSE); 
    and SMC_I5(ENABLE_E_AND_NOT_SE,dE, SE_bar); 
 
    not SMC_I6(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I7(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDQHDV2 ( Q, CK, D, E, SE, SI, VDD, VSS); 
input CK, D, E, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_sedff_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I4(SE_bar,dSE); 
    and SMC_I5(ENABLE_E_AND_NOT_SE,dE, SE_bar); 
 
    not SMC_I6(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I7(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDQHDV4 ( Q, CK, D, E, SE, SI, VDD, VSS); 
input CK, D, E, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_sedff_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I4(SE_bar,dSE); 
    and SMC_I5(ENABLE_E_AND_NOT_SE,dE, SE_bar); 
 
    not SMC_I6(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I7(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDQHDV8 ( Q, CK, D, E, SE, SI, VDD, VSS); 
input CK, D, E, SE, SI;
inout VDD, VSS;
output Q;
wire Q_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  udp_sedff_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  buf     I1 (Q_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I4(SE_bar,dSE); 
    and SMC_I5(ENABLE_E_AND_NOT_SE,dE, SE_bar); 
 
    not SMC_I6(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I7(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CK --> Q 
	(posedge CK => (Q : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDQNHDV0 ( QN, CK, D, E, SE, SI, VDD, VSS); 
input CK, D, E, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN; 
  udp_sedff_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I6(SE_bar,dSE); 
    and SMC_I7(ENABLE_E_AND_NOT_SE,dE, SE_bar); 
 
    not SMC_I8(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I9(ENABLE_SE,dSE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDQNHDV2 ( QN, CK, D, E, SE, SI, VDD, VSS); 
input CK, D, E, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN; 
  udp_sedff_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I6(SE_bar,dSE); 
    and SMC_I7(ENABLE_E_AND_NOT_SE,dE, SE_bar); 
 
    not SMC_I8(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I9(ENABLE_SE,dSE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDQNHDV4 ( QN, CK, D, E, SE, SI, VDD, VSS); 
input CK, D, E, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN; 
  udp_sedff_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I6(SE_bar,dSE); 
    and SMC_I7(ENABLE_E_AND_NOT_SE,dE, SE_bar); 
 
    not SMC_I8(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I9(ENABLE_SE,dSE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDQNHDV8 ( QN, CK, D, E, SE, SI, VDD, VSS); 
input CK, D, E, SE, SI;
inout VDD, VSS;
output QN;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN; 
  udp_sedff_PWR I0 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  not     I2 (QN_temp, n0 );
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I6(SE_bar,dSE); 
    and SMC_I7(ENABLE_E_AND_NOT_SE,dE, SE_bar); 
 
    not SMC_I8(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I9(ENABLE_SE,dSE); 
 
 
  specify 
 
 
 
	// arc CK --> QN 
	(posedge CK => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CK,1.0,0,NOTIFIER); 
 
        $width(posedge CK,1.0,0,NOTIFIER); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
        $setuphold(posedge CK &&& (ENABLE_E_AND_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_E_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dD); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            negedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
        $setuphold(posedge CK &&& (ENABLE_NOT_SE === 1'b1), 
            posedge E &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dE); 
 
 
 
        $setuphold(posedge CK, negedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
        $setuphold(posedge CK, posedge SE, 1.0, 1.0, NOTIFIER, , , dCK, dSE); 
 
 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
        $setuphold(posedge CK &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCK, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDRNQHDV0 (D, E, RDN, SE, SI, CK, Q, VDD, VSS); 
  input D, E, RDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI;
  buf       I0 (xRN, dRDN );
  udp_sedff_PWR I1 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  buf       I2 (Q_temp, n0 );
  assign ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI=(D&E&!SE|E&SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_E_AND_RDN_AND_NOT_SE,dE,dRDN, SE_bar);

    and SMC_I6(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I7(ENABLE_RDN,dRDN);

    and SMC_I8(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDRNQHDV2 (D, E, RDN, SE, SI, CK, Q, VDD, VSS); 
  input D, E, RDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI;
  buf       I0 (xRN, dRDN );
  udp_sedff_PWR I1 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  buf       I2 (Q_temp, n0 );
  assign ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI=(D&E&!SE|E&SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_E_AND_RDN_AND_NOT_SE,dE,dRDN, SE_bar);

    and SMC_I6(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I7(ENABLE_RDN,dRDN);

    and SMC_I8(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDRNQHDV4 (D, E, RDN, SE, SI, CK, Q, VDD, VSS); 
  input D, E, RDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI;
  buf       I0 (xRN, dRDN );
  udp_sedff_PWR I1 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  buf       I2 (Q_temp, n0 );
  assign ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI=(D&E&!SE|E&SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_E_AND_RDN_AND_NOT_SE,dE,dRDN, SE_bar);

    and SMC_I6(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I7(ENABLE_RDN,dRDN);

    and SMC_I8(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDRNQHDV8 (D, E, RDN, SE, SI, CK, Q, VDD, VSS); 
  input D, E, RDN, SE, SI, CK;

inout VDD, VSS;
  output Q;
wire Q_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI;
  buf       I0 (xRN, dRDN );
  udp_sedff_PWR I1 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
  buf       I2 (Q_temp, n0 );
  assign ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI=(D&E&!SE|E&SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar,dSE);
    and SMC_I5(ENABLE_E_AND_RDN_AND_NOT_SE,dE,dRDN, SE_bar);

    and SMC_I6(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I7(ENABLE_RDN,dRDN);

    and SMC_I8(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CK --> Q
	(posedge CK => (Q : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDRNQNHDV0 (D, E, RDN, SE, SI, CK, QN, VDD, VSS); 
  input D, E, RDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  wire ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI;
   buf       I0 (xRN, dRDN );
   udp_sedff_PWR I1 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
   not       I3 (QN_temp, n0 );
   assign ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI=(D&E&!SE|E&SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_E_AND_RDN_AND_NOT_SE,dE,dRDN, SE_bar);

    and SMC_I8(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I9(ENABLE_RDN,dRDN);

    and SMC_I10(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDRNQNHDV2 (D, E, RDN, SE, SI, CK, QN, VDD, VSS); 
  input D, E, RDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  wire ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI;
   buf       I0 (xRN, dRDN );
   udp_sedff_PWR I1 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
   not       I3 (QN_temp, n0 );
   assign ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI=(D&E&!SE|E&SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_E_AND_RDN_AND_NOT_SE,dE,dRDN, SE_bar);

    and SMC_I8(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I9(ENABLE_RDN,dRDN);

    and SMC_I10(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDRNQNHDV4 (D, E, RDN, SE, SI, CK, QN, VDD, VSS); 
  input D, E, RDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  wire ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI;
   buf       I0 (xRN, dRDN );
   udp_sedff_PWR I1 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
   not       I3 (QN_temp, n0 );
   assign ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI=(D&E&!SE|E&SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_E_AND_RDN_AND_NOT_SE,dE,dRDN, SE_bar);

    and SMC_I8(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I9(ENABLE_RDN,dRDN);

    and SMC_I10(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SEDRNQNHDV8 (D, E, RDN, SE, SI, CK, QN, VDD, VSS); 
  input D, E, RDN, SE, SI, CK;

inout VDD, VSS;
  output QN;
wire QN_temp;

  reg NOTIFIER;
  wire ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI;
   buf       I0 (xRN, dRDN );
   udp_sedff_PWR I1 (n0, dD, dCK, xRN, dSI, dSE, dE, VDD, VSS, NOTIFIER ); 
   not       I3 (QN_temp, n0 );
   assign ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI=(D&E&!SE|E&SE&SI)? 1'b1:1'b0;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar,dSE);
    and SMC_I7(ENABLE_E_AND_RDN_AND_NOT_SE,dE,dRDN, SE_bar);

    and SMC_I8(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I9(ENABLE_RDN,dRDN);

    and SMC_I10(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify



	// arc CK --> QN
	(posedge CK => (QN : D))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b0 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b0 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CK===1'b1 && D===1'b1 && E===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CK,1.0,0,NOTIFIER);

        $width(posedge CK,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);

        $setuphold(posedge CK &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_E_AND_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dD);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge E &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dE);



        $setuphold(posedge CK &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_E_AND_NOT_SE_OR_E_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCK, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);

        $setuphold(posedge CK &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSE);



        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);

        $setuphold(posedge CK &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCK, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDHDV0 ( Q, QN, CKN, D, SE, SI, VDD, VSS); 
input CKN, D, SE, SI;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I7(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I8(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CKN --> Q 
	(negedge CKN => (Q : D))  = (1.0,1.0); 
 
	// arc CKN --> QN 
	(negedge CKN => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CKN,1.0,0,NOTIFIER); 
 
        $width(posedge CKN,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CKN &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dD); 
 
        $setuphold(negedge CKN &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dD); 
 
 
 
        $setuphold(negedge CKN, negedge SE, 1.0, 1.0, NOTIFIER, , , dCKN, dSE); 
 
        $setuphold(negedge CKN, posedge SE, 1.0, 1.0, NOTIFIER, , , dCKN, dSE); 
 
 
 
        $setuphold(negedge CKN &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dSI); 
 
        $setuphold(negedge CKN &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDHDV2 ( Q, QN, CKN, D, SE, SI, VDD, VSS); 
input CKN, D, SE, SI;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I7(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I8(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CKN --> Q 
	(negedge CKN => (Q : D))  = (1.0,1.0); 
 
	// arc CKN --> QN 
	(negedge CKN => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CKN,1.0,0,NOTIFIER); 
 
        $width(posedge CKN,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CKN &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dD); 
 
        $setuphold(negedge CKN &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dD); 
 
 
 
        $setuphold(negedge CKN, negedge SE, 1.0, 1.0, NOTIFIER, , , dCKN, dSE); 
 
        $setuphold(negedge CKN, posedge SE, 1.0, 1.0, NOTIFIER, , , dCKN, dSE); 
 
 
 
        $setuphold(negedge CKN &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dSI); 
 
        $setuphold(negedge CKN &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDHDV4 ( Q, QN, CKN, D, SE, SI, VDD, VSS); 
input CKN, D, SE, SI;
inout VDD, VSS;
output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER; 
  supply1 xRN, xSN; 
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional // 
 
  `else // functional // 
    not SMC_I7(ENABLE_NOT_SE,dSE); 
 
    buf SMC_I8(ENABLE_SE,dSE); 
 
 
  specify 
 
 
	// arc CKN --> Q 
	(negedge CKN => (Q : D))  = (1.0,1.0); 
 
	// arc CKN --> QN 
	(negedge CKN => (QN : D))  = (1.0,1.0); 
 
        $width(negedge CKN,1.0,0,NOTIFIER); 
 
        $width(posedge CKN,1.0,0,NOTIFIER); 
 
        $setuphold(negedge CKN &&& (ENABLE_NOT_SE === 1'b1), 
            negedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dD); 
 
        $setuphold(negedge CKN &&& (ENABLE_NOT_SE === 1'b1), 
            posedge D &&& (ENABLE_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dD); 
 
 
 
        $setuphold(negedge CKN, negedge SE, 1.0, 1.0, NOTIFIER, , , dCKN, dSE); 
 
        $setuphold(negedge CKN, posedge SE, 1.0, 1.0, NOTIFIER, , , dCKN, dSE); 
 
 
 
        $setuphold(negedge CKN &&& (ENABLE_SE === 1'b1), 
            negedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dSI); 
 
        $setuphold(negedge CKN &&& (ENABLE_SE === 1'b1), 
            posedge SI &&& (ENABLE_SE === 1'b1), 1.0, 1.0, NOTIFIER, , , 
            dCKN, dSI); 
 
 
 
 
  endspecify 
 
  `endif // functional // 
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDRNHDV0 (D, RDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);
    and SMC_I8(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I9(ENABLE_RDN,dRDN);

    and SMC_I10(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDRNHDV2 (D, RDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);
    and SMC_I8(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I9(ENABLE_RDN,dRDN);

    and SMC_I10(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDRNHDV4 (D, RDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xSN;
wire ENABLE_D_AND_NOT_SE_OR_SE_AND_SI;
  buf   XX0 (xRN, dRDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_NOT_SE_OR_SE_AND_SI=(D&!SE | SE&SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);
    and SMC_I8(ENABLE_RDN_AND_NOT_SE,dRDN, SE_bar);

    buf SMC_I9(ENABLE_RDN,dRDN);

    and SMC_I10(ENABLE_RDN_AND_SE,dRDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), posedge RDN &&& (ENABLE_D_AND_NOT_SE_OR_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            negedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_RDN === 1'b1),
            posedge SE &&& (ENABLE_RDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDRSNHDV0 (D, RDN, SDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(SE_bar,dSE);

    and SMC_I9(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I10(ENABLE_SDN,dSDN);

    buf SMC_I11(ENABLE_RDN,dRDN);

    and SMC_I12(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I13(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDRSNHDV2 (D, RDN, SDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(SE_bar,dSE);

    and SMC_I9(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I10(ENABLE_SDN,dSDN);

    buf SMC_I11(ENABLE_RDN,dRDN);

    and SMC_I12(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I13(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDRSNHDV4 (D, RDN, SDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, RDN, SDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
wire ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI;
wire ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI;
  buf   XX0 (xRN, dRDN );
  buf   XX1 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI=(D&SDN&!SE|SDN&SE&SI)? 1'b1:1'b0;
  assign ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI=(!D&RDN&!SE|RDN&SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(SE_bar,dSE);

    and SMC_I9(ENABLE_RDN_AND_SDN_AND_NOT_SE,dRDN,dSDN, SE_bar);

    buf SMC_I10(ENABLE_SDN,dSDN);

    buf SMC_I11(ENABLE_RDN,dRDN);

    and SMC_I12(ENABLE_RDN_AND_SDN,dRDN,dSDN);

    and SMC_I13(ENABLE_RDN_AND_SDN_AND_SE,dRDN,dSDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> Q
	(negedge RDN => (Q : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc RDN --> QN
	(negedge RDN => (QN : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && RDN===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_RDN_AND_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1),
            posedge RDN &&& (ENABLE_D_AND_SDN_AND_NOT_SE_OR_SDN_AND_SE_AND_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dRDN);


        $width(negedge RDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1),
            posedge SDN &&& (ENABLE_NOT_D_AND_RDN_AND_NOT_SE_OR_RDN_AND_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSDN);


        $setuphold(posedge RDN, posedge SDN, 1.0, 1.0, NOTIFIER, , , dRDN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            negedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN === 1'b1),
            posedge SE &&& (ENABLE_RDN_AND_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_RDN_AND_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDSNHDV0 (D, SDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, SDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);
    and SMC_I8(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    and SMC_I10(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDSNHDV2 (D, SDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, SDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);
    and SMC_I8(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    and SMC_I10(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
/*****************************************************************************/
`timescale 10 ps / 1 ps

`ifdef functional
                                // none
`else
        `define SMC_NFORCE 1    // Flag to force output to x if notifer changes
`endif

`celldefine 
module SNDSNHDV4 (D, SDN, SE, SI, CKN, Q, QN, VDD, VSS); 
  input D, SDN, SE, SI, CKN;

inout VDD, VSS;
  output Q, QN;
wire Q_temp;
wire QN_temp;

  reg NOTIFIER;
  supply1 xRN;
wire ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI;
  buf   XX0 (xSN, dSDN );
  not     IC (clk, dCKN );
  udp_dff_PWR I0 (n0, n1, clk, xRN, xSN, VDD, VSS, NOTIFIER ); 
  udp_mux_PWR I1 (n1, dD, dSI, dSE ,VDD, VSS); 
  buf     I2 (Q_temp, n0 );
  not     I3 (QN_temp, n0 );
  assign ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI=(!D&!SE|SE&!SI)? 1'b1:1'b0;
  assign Q = ((VDD === 1'b1) && (VSS === 1'b0)) ? Q_temp : 1'bx;
  assign QN = ((VDD === 1'b1) && (VSS === 1'b0)) ? QN_temp : 1'bx;
  `ifdef functional // functional //

  `else // functional //
    not SMC_I7(SE_bar,dSE);
    and SMC_I8(ENABLE_SDN_AND_NOT_SE,dSDN, SE_bar);

    buf SMC_I9(ENABLE_SDN,dSDN);

    and SMC_I10(ENABLE_SDN_AND_SE,dSDN,dSE);


  specify


	// arc CKN --> Q
	(negedge CKN => (Q : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> Q
	(negedge SDN => (Q : 1'b1))  = (1.0,1.0);

	// arc CKN --> QN
	(negedge CKN => (QN : D))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b0 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b0 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b0 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b0)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

	if(CKN===1'b1 && D===1'b1 && SE===1'b1 && SI===1'b1)
	// arc SDN --> QN
	(negedge SDN => (QN : 1'b0))  = (1.0,1.0);

        $width(negedge CKN,1.0,0,NOTIFIER);

        $width(posedge CKN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            negedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_NOT_SE === 1'b1),
            posedge D &&& (ENABLE_SDN_AND_NOT_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dD);



        $setuphold(negedge CKN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), posedge SDN &&& (ENABLE_NOT_D_AND_NOT_SE_OR_SE_AND_NOT_SI === 1'b1), 1.0, 1.0, NOTIFIER, , , dCKN, dSDN);


        $width(negedge SDN,1.0,0,NOTIFIER);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            negedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);

        $setuphold(negedge CKN &&& (ENABLE_SDN === 1'b1),
            posedge SE &&& (ENABLE_SDN === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSE);



        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_SE === 1'b1),
            negedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);

        $setuphold(negedge CKN &&& (ENABLE_SDN_AND_SE === 1'b1),
            posedge SI &&& (ENABLE_SDN_AND_SE === 1'b1), 1.0, 1.0, NOTIFIER, , ,
            dCKN, dSI);




  endspecify

  `endif // functional //
endmodule
`endcelldefine
// $Id: udp_dff.v
// verilog UDP for d flip-flops 
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//
primitive udp_dff_PWR (out, in, clk, clr_, set_, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, VDD, VSS, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  VDD  VSS  NOT  : Qt : Qt+1
//
   0  r   ?   1   1	0	?   : ?  :  0  ; // clock in 0
   1  r   1   ?   1	0	?   : ?  :  1  ; // clock in 1
   1  *   1   ?   1	0	?   : 1  :  1  ; // reduce pessimism
   0  *   ?   1   1	0	?   : 0  :  0  ; // reduce pessimism
   ?  f   ?   ?   1	0	?   : ?  :  -  ; // no changes on negedge clk
   *  b   ?   ?   1	0	?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   0   1	0	?   : ?  :  1  ; // set output
   ?  b   1   *   1	0	?   : 1  :  1  ; // cover all transistions on set_
   1  x   1   *   1	0	?   : 1  :  1  ; // cover all transistions on set_
   ?  ?   0   1   1	0	?   : ?  :  0  ; // reset output
   ?  b   *   1   1	0	?   : 0  :  0  ; // cover all transistions on clr_
   0  x   *   1   1	0	?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?   ?   ?   0	0	?   : ?  :  x  ;
   ?  ?   ?   ?   0	1	?   : ?  :  x  ;
   ?  ?   ?   ?   1	1	?   : ?  :  x  ;
   ?  ?   ?   ?   ?	?	*   : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_dff

primitive udp_dff_rdn_pre_sdn_PWR (out, in, clk, clr_, set_, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, VDD, VSS, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  VDD  VSS  NOT  : Qt : Qt+1
//
   0  r   ?   1   1	0	?   : ?  :  0  ; // clock in 0
   1  r   1   ?   1	0	?   : ?  :  1  ; // clock in 1
   1  *   1   ?   1	0	?   : 1  :  1  ; // reduce pessimism
   0  *   ?   1   1	0	?   : 0  :  0  ; // reduce pessimism
   ?  f   ?   ?   1	0	?   : ?  :  -  ; // no changes on negedge clk
   *  b   ?   ?   1	0 	?   : ?  :  -  ; // no changes when in switches
   ?  ?   1   0   1	0 	?   : ?  :  1  ; // set output
   ?  b   1   *   1	0	?   : 1  :  1  ; // cover all transistions on set_
   1  x   1   *   1	0	?   : 1  :  1  ; // cover all transistions on set_
   ?  ?   0   ?   1	0 	?   : ?  :  0  ; // reset output
   ?  b   *   1   1	0 	?   : 0  :  0  ; // cover all transistions on clr_
   0  x   *   1   1	0	?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?   ?   ?   0	0	?   : ?  :  x  ;
   ?  ?   ?   ?   0	1	?   : ?  :  x  ;
   ?  ?   ?   ?   1	1	?   : ?  :  x  ;
   ?  ?   ?   ?   ?	?	*   : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_dff_rdn_pre_sdn


// $Id: udp_edff.v
// verilog UDP for d flip-flops with enable
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_edff_PWR (out, in, clk, clr_, set_, en, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, en, VDD, VSS, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  en  VDD VSS NOT  : Qt : Qt+1
//
   0   r    ?      1     1   1	0	?    : ?  :  0  ; // clock in 0
   1   r    1      ?     1   1	0	?    : ?  :  1  ; // clock in 1
   ?   *    1      ?     0   1	0	?    : ?  :  -  ; // no changes, not enabled
   *   ?    1      ?     0   1	0	?    : ?  :  -  ; // no changes, not enabled
   1   *    1      ?     ?   1	0	?    : 1  :  1  ; // reduce pessimism
   0   *    ?      1     ?   1	0	?    : 0  :  0  ; // reduce pessimism
   ?   f    ?      ?     ?   1	0	?    : ?  :  -  ; // no changes on negedge clk
   *   b    ?      ?     ?   1	0	?    : ?  :  -  ; // no changes when in switches
   1   x    1      ?     ?   1	0	?    : 1  :  1  ; // no changes when in switches
   0   x    ?      1     ?   1	0	?    : 0  :  0  ; // no changes when in switches
   ?   b    ?      ?     *   1	0	?    : ?  :  -  ; // no changes when en switches
   ?   x    1      1     0   1	0	?    : ?  :  -  ; // no changes when en is disabled
   ?   ?    ?      0     ?   1	0	?    : ?  :  1  ; // set output
   ?   b    1      *     ?   1	0	?    : 1  :  1  ; // cover all transistions on set_
   ?   ?    1      *     0   1	0	?    : 1  :  1  ; // cover all transistions on set_
   ?   ?    0      1     ?   1	0	?    : ?  :  0  ; // reset output
   ?   b    *      1     ?   1	0	?    : 0  :  0  ; // cover all transistions on clr_
   ?   ?    *      1     0   1	0	?    : 0  :  0  ; // cover all transistions on clr_
   ?   ?    ?      ?     ?   0	0	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   0	1	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   1	1	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   ?	?	*    : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_edff

// $Id: udp_edfft.v
// verilog UDP for d flip-flops with enable
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_edfft_PWR (out, in, clk, clr_, set_, en, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, en, VDD, VSS, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  en  VDD VSS NOT  : Qt : Qt+1
//
   ?   r    0      1     ?   1	0	?    : ?  :  0  ; // clock in 0
   0   r    ?      1     1   1	0	?    : ?  :  0  ; // clock in 0
   ?   r    ?      0     ?   1	0	?    : ?  :  1  ; // clock in 1
   1   r    1      ?     1   1	0	?    : ?  :  1  ; // clock in 1
   ?   *    1      1     0   1	0	?    : ?  :  -  ; // no changes, not enabled
   ?   *    ?      1     0   1	0	?    : 0  :  0  ; // no changes, not enabled
   ?   *    1      ?     0   1	0	?    : 1  :  1  ; // no changes, not enabled
   ?  (x0)  ?      ?     ?   1	0	?    : ?  :  -  ; // no changes
   ?  (x1)  ?      0     ?   1	0	?    : 1  :  1  ; // no changes
   1   *    1      ?     ?   1	0	?    : 1  :  1  ; // reduce pessimism
   0   *    ?      1     ?   1	0	?    : 0  :  0  ; // reduce pessimism
   ?   f    ?      ?     ?   1	0	?    : ?  :  -  ; // no changes on negedge clk
   *   b    ?      ?     ?   1	0	?    : ?  :  -  ; // no changes when in switches
   1   x    1      ?     ?   1	0	?    : 1  :  1  ; // no changes when in switches
   ?   x    1      ?     0   1	0	?    : 1  :  1  ; // no changes when in switches
   0   x    ?      1     ?   1	0	?    : 0  :  0  ; // no changes when in switches
   ?   x    ?      1     0   1	0	?    : 0  :  0  ; // no changes when in switches
   ?   b    ?      ?     *   1	0	?    : ?  :  -  ; // no changes when en switches
   ?   b    *      ?     ?   1	0	?    : ?  :  -  ; // no changes when clr_ switches
   ?   x    0      1     ?   1	0	?    : 0  :  0  ; // no changes when clr_ switches
   ?   b    ?      *     ?   1	0	?    : ?  :  -  ; // no changes when set_ switches
   ?   x    ?      0     ?   1	0	?    : 1  :  1  ; // no changes when set_ switches
   ?   ?    ?      ?     ?   0	0	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   0	1	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   1	1	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   ?	?	*    : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_edfft

// $Id: udp_edffts.v
//
// verilog UDP for d flip-flops with enable
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_edffts_PWR (out, in, clk, clr_, set_, en, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, en, VDD, VSS, NOTIFIER;
   reg    out;

   table

// in  clk  clr_   set_  en  VDD VSS NOT  : Qt : Qt+1
//
   ?   r    0      ?     ?   1	0	?    : ?  :  0  ; // clock in 0
   0   r    ?      1     1   1	0	?    : ?  :  0  ; // clock in 0
   ?   r    1      0     ?   1	0	?    : ?  :  1  ; // clock in 1
   1   r    1      ?     1   1	0	?    : ?  :  1  ; // clock in 1
   ?   *    1      1     0   1	0	?    : ?  :  -  ; // no changes, not enabled
   ?   *    ?      1     0   1	0	?    : 0  :  0  ; // no changes, not enabled
   ?   *    1      ?     0   1	0	?    : 1  :  1  ; // no changes, not enabled
   ?  (x0)  ?      ?     ?   1	0	?    : ?  :  -  ; // no changes
   ?  (x1)  ?      0     ?   1	0	?    : 1  :  1  ; // no changes
   1   *    1      ?     ?   1	0	?    : 1  :  1  ; // reduce pessimism
   0   *    ?      1     ?   1	0	?    : 0  :  0  ; // reduce pessimism
   ?   f    ?      ?     ?   1	0	?    : ?  :  -  ; // no changes on negedge clk
   *   b    ?      ?     ?   1	0	?    : ?  :  -  ; // no changes when in switches
   1   x    1      ?     ?   1	0	?    : 1  :  1  ; // no changes when in switches
   ?   x    1      ?     0   1	0	?    : 1  :  1  ; // no changes when in switches
   0   x    ?      1     ?   1	0	?    : 0  :  0  ; // no changes when in switches
   ?   x    ?      1     0   1	0	?    : 0  :  0  ; // no changes when in switches
   ?   b    ?      ?     *   1	0	?    : ?  :  -  ; // no changes when en switches
   ?   b    *      ?     ?   1	0	?    : ?  :  -  ; // no changes when clr_ switches
   ?   x    0      1     ?   1	0	?    : 0  :  0  ; // no changes when clr_ switches
   ?   b    ?      *     ?   1	0	?    : ?  :  -  ; // no changes when set_ switches
   ?   x    ?      0     ?   1	0	?    : 1  :  1  ; // no changes when set_ switches
   ?   ?    ?      ?     ?   0	1	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   0	0	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   1	1	?    : ?  :  x  ;
   ?   ?    ?      ?     ?   ?	?	*    : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_edffts

// $Id: udp_jkff.v
//
// verilog UDP for jk flip-flps
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_jkff_PWR (out, j, k, clk, clr_, set_, VDD, VSS, NOTIFIER);
   output out;  
   input  j, k, clk, clr_, set_, VDD, VSS, NOTIFIER;
   reg    out;

   table

// j  k  clk  clr_   set_  VDD  VSS  NOT  : Qt : Qt+1
//       
   0  0  r   1   1   1	0	?   : ?  :  -  ; // output remains same
   0  1  r   ?   1   1	0	?   : ?  :  0  ; // clock in 0
   1  0  r   1   ?   1	0	?   : ?  :  1  ; // clock in 1
   ?  1  r   ?   1   1	0	?   : 1  :  0  ; // clock in 0
   1  ?  r   1   ?   1	0	?   : 0  :  1  ; // clock in 1
   ?  0  *   1   ?   1	0	?   : 1  :  1  ; // reduce pessimism
   0  ?  *   ?   1   1	0	?   : 0  :  0  ; // reduce pessimism
   ?  ?  f   ?   ?   1	0	?   : ?  :  -  ; // no changes on negedge clk
   *  ?  b   ?   ?   1	0	?   : ?  :  -  ; // no changes when j switches
   *  0  x   1   ?   1	0	?   : 1  :  1  ; // no changes when j switches
   ?  *  b   ?   ?   1	0	?   : ?  :  -  ; // no changes when k switches
   0  *  x   ?   1   1	0	?   : 0  :  0  ; // no changes when k switches
   ?  ?  ?   ?   0   1	0	?   : ?  :  1  ; // set output
   ?  ?  b   1   *   1	0	?   : 1  :  1  ; // cover all transistions on set_
   ?  0  x   1   *   1	0	?   : 1  :  1  ; // cover all transistions on set_
   ?  ?  ?   0   1   1	0	?   : ?  :  0  ; // reset output
   ?  ?  b   *   1   1	0	?   : 0  :  0  ; // cover all transistions on clr_
   0  ?  x   *   1   1	0	?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?  ?   ?   ?   0	1	?   : ?  :  x  ;
   ?  ?  ?   ?   ?   1	1	?   : ?  :  x  ;
   ?  ?  ?   ?   ?   0	0	?   : ?  :  x  ;
   ?  ?  ?   ?   ?   ?	?	*   : ?  :  x  ; // any NOTIFIER change

   endtable
endprimitive // udp_jkff

// $Id: udp_sedff.v
//
// verilog UDP for a 2-input mux used in scan cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//
 primitive udp_sedff_PWR (out, in, clk, clr_, si, se, en, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, clr_, si, se,  en, VDD, VSS, NOTIFIER;
   reg    out;

   table
   // in  clk  clr_  si  se  en  VDD  VSS  NOT : Qt : Qt+1
      ?    ?    ?     ?   ?   ?   ?	?   *  : ?  :  x; // any NOTIFIER changed
      ?    ?    0     ?   ?   ?   1     0   ?  : ?  :  0;     
      ?    r    ?     0   1   ?   1     0   ?  : ?  :  0;     
      ?    r    1     1   1   ?   1     0   ?  : ?  :  1;
      ?    b    1     ?   *   ?   1     0   ?  : ?  :  -; // no changes when se switches
      ?    b    1     *   ?   ?   1     0   ?  : ?  :  -; // no changes when si switches
      *    b    1     ?   ?   ?   1     0   ?  : ?  :  -; // no changes when in switches
      *    ?    ?     ?   0   0   1     0   ?  : 0  :  0; // no changes when in switches
      ?    ?    ?     *   0   0   1     0   ?  : 0  :  0; // no changes when in switches
      ?    b    1     ?   ?   *   1     0   ?  : ?  :  -; // no changes when en switches
      ?    b    *     ?   ?   ?   1     0   ?  : 0  :  0; // no changes when en switches
      ?    ?    *     ?   0   0   1     0   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     ?   ?   *   1     0   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     ?   *   ?   1     0   ?  : 0  :  0; // no changes when en switches
      ?    b    ?     *   ?   ?   1     0   ?  : 0  :  0; // no changes when en switches
      *    b    ?     ?   ?   ?   1     0   ?  : 0  :  0; // no changes when en switches
      ?  (10)   ?     ?   ?   ?   1     0   ?  : ?  :  -;  // no changes on falling clk edge
      ?    *    1     1   1   ?   1     0   ?  : 1  :  1;
      ?    x    1     1   1   ?   1     0   ?  : 1  :  1;
      ?    *    1     1   ?   0   1     0   ?  : 1  :  1;
      ?    x    1     1   ?   0   1     0   ?  : 1  :  1;
      ?    *    ?     0   1   ?   1     0   ?  : 0  :  0;
      ?    x    ?     0   1   ?   1     0   ?  : 0  :  0;
      ?    *    ?     0   ?   0   1     0   ?  : 0  :  0;
      ?    x    ?     0   ?   0   1     0   ?  : 0  :  0;
      0    r    ?     0   ?   1   1     0   ?  : ?  :  0 ; 
      0    *    ?     0   ?   ?   1     0   ?  : 0  :  0 ; 
      0    x    ?     0   ?   ?   1     0   ?  : 0  :  0 ; 
      1    r    1     1   ?   1   1     0   ?  : ?  :  1 ; 
      1    *    1     1   ?   ?   1     0   ?  : 1  :  1 ; 
      1    x    1     1   ?   ?   1     0   ?  : 1  :  1 ; 
      ?  (x0)   ?     ?   ?   ?   1     0   ?  : ?  :  -;  // no changes on falling clk edge
      1    r    1     ?   0   1   1     0   ?  : ?  :  1;
      0    r    ?     ?   0   1   1     0   ?  : ?  :  0;
      ?    *    ?     ?   0   0   1     0   ?  : ?  :  -;
      ?    x    1     ?   0   0   1     0   ?  : ?  :  -;
      1    x    1     ?   0   ?   1     0   ?  : 1  :  1; // no changes when in switches
      0    x    ?     ?   0   ?   1     0   ?  : 0  :  0; // no changes when in switches
      1    x    ?     ?   0   0   1     0   ?  : 0  :  0; // no changes when in switches
      1    *    1     ?   0   ?   1     0   ?  : 1  :  1; // reduce pessimism
      0    *    ?     ?   0   ?   1     0   ?  : 0  :  0; // reduce pessimism
      ?    ?    ?     ?   ?   ?   0	1   ?  : ?  :  x;
      ?    ?    ?     ?   ?   ?   1	1   ?  : ?  :  x;
      ?    ?    ?     ?   ?   ?   0	0   ?  : ?  :  x;

   endtable
endprimitive  /* udp_sedff */
   
// $Id: udp_sedfft.v
//
// verilog UDP for a 2-input mux used in scan cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//
 primitive udp_sedfft_PWR (out, in, clk, clr_, si, se, en, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, clr_, si, se,  en, VDD, VSS, NOTIFIER;
   reg    out;

   table
   // in  clk  clr_  si  se  en  VDD  VSS  NOT : Qt : Qt+1
      ?    ?    ?     ?   ?   ?   ?    ?    *  : ?  :  x; // any NOTIFIER changed
      ?    r    ?     0   1   ?   1    0    ?  : ?  :  0;     
      ?    r    ?     1   1   ?   1    0    ?  : ?  :  1;
      ?    b    ?     ?   *   ?   1    0    ?  : ?  :  -; // no changes when se switches
      ?    b    ?     *   ?   ?   1    0    ?  : ?  :  -; // no changes when si switches
      *    b    ?     ?   ?   ?   1    0    ?  : ?  :  -; // no changes when in switches
      ?    b    ?     ?   ?   *   1    0    ?  : ?  :  -; // no changes when en switches
      ?    b    *     ?   ?   ?   1    0    ?  : ?  :  -; // no changes when clr switches
      0    r    ?     0   ?   1   1    0    ?  : ?  :  0 ; 
      1    r    1     1   ?   1   1    0    ?  : ?  :  1 ; 
      ?    r    ?     0   ?   0   1    0    ?  : 0  :  0;
      ?    x    ?     0   ?   0   1    0    ?  : 0  :  0;
      ?    r    1     1   ?   0   1    0    ?  : 1  :  1;
      ?    x    1     1   ?   0   1    0    ?  : 1  :  1;
      ?    *    1     ?   0   0   1    0    ?  : ?  :  -;
      ?    *    ?     1   1   ?   1    0    ?  : 1  :  1;
      1    *    1     1   ?   ?   1    0    ?  : 1  :  1;
      ?    *    ?     0   1   ?   1    0    ?  : 0  :  0;
      ?    *    0     0   ?   ?   1    0    ?  : 0  :  0;
      0    *    ?     0   ?   ?   1    0    ?  : 0  :  0;
      ?    x    1     ?   0   0   1    0    ?  : ?  :  -;
      ?    *    ?     ?   0   0   1    0    ?  : 0  :  0;
      ?    x    ?     ?   0   0   1    0    ?  : 0  :  0;
      ?    x    ?     1   1   ?   1    0    ?  : 1  :  1;
      1    x    1     1   ?   ?   1    0    ?  : 1  :  1;
      ?    x    ?     0   1   ?   1    0    ?  : 0  :  0;
      ?    x    0     0   ?   ?   1    0    ?  : 0  :  0;
      0    x    ?     0   ?   ?   1    0    ?  : 0  :  0;
      ?    r    0     0   ?   ?   1    0    ?  : ?  :  0 ; 
      ?   (?0)  ?     ?   ?   ?   1    0    ?  : ?  :  -;  // no changes on falling clk edge
      1    r    1     ?   0   1   1    0    ?  : ?  :  1;
      0    r    ?     ?   0   1   1    0    ?  : ?  :  0;
      ?    r    0     ?   0   ?   1    0    ?  : ?  :  0;
      ?    x    0     ?   0   ?   1    0    ?  : 0  :  0;
      1    x    1     ?   0   ?   1    0    ?  : 1  :  1; // no changes when in switches
      0    x    ?     ?   0   ?   1    0    ?  : 0  :  0; // no changes when in switches
      1    *    1     ?   0   ?   1    0    ?  : 1  :  1; // reduce pessimism
      0    *    ?     ?   0   ?   1    0    ?  : 0  :  0; // reduce pessimism
      ?    ?    ?     ?   ?   ?   0    1    ?  : ?  :  x;
      ?    ?    ?     ?   ?   ?   1    1    ?  : ?  :  x;
      ?    ?    ?     ?   ?   ?   0    0    ?  : ?  :  x;

   endtable
endprimitive  /* udp_sedfft */

/*   
// $Id: udp_sedffts.v
//
// verilog UDP for a 2-input mux used in scan cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//
 primitive udp_sedffts_PWR (out, in, clk, set_, si, se, en, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, set_, si, se,  en, VDD, VSS, NOTIFIER;
   reg    out;

   table
   // in  clk  set_  si  se  en  VDD  VSS  NOT : Qt : Qt+1
      ?    ?    ?     ?   ?   ?   ?    ?    *  : ?  :  x; // any NOTIFIER changed
      ?    r    ?     0   1   ?   1    0    ?  : ?  :  0;     
      ?    r    ?     1   1   ?   1    0    ?  : ?  :  1;
      ?    b    ?     ?   *   ?   1    0    ?  : ?  :  -; // no changes when se switches
      ?    b    ?     *   ?   ?   1    0    ?  : ?  :  -; // no changes when si switches
      *    b    ?     ?   ?   ?   1    0    ?  : ?  :  -; // no changes when in switches
      ?    b    ?     ?   ?   *   1    0    ?  : ?  :  -; // no changes when en switches
      ?    b    *     ?   ?   ?   1    0    ?  : ?  :  -; // no changes when clr switches
      0    r    ?     0   ?   1   1    0    ?  : ?  :  0 ; 
      1    r    1     1   ?   1   1    0    ?  : ?  :  1 ; 
      ?    r    ?     0   ?   0   1    0    ?  : 0  :  0;
      ?    x    ?     0   ?   0   1    0    ?  : 0  :  0;
      ?    r    1     1   ?   0   1    0    ?  : 1  :  1;
      ?    x    1     1   ?   0   1    0    ?  : 1  :  1;
      ?    *    1     ?   0   0   1    0    ?  : ?  :  -;
      ?    *    ?     1   1   ?   1    0    ?  : 1  :  1;
      1    *    1     1   ?   ?   1    0    ?  : 1  :  1;
      ?    *    ?     0   1   ?   1    0    ?  : 0  :  0;
      ?    *    0     0   ?   ?   1    0    ?  : 0  :  1;
      0    *    ?     0   ?   ?   1    0    ?  : 0  :  0;
      ?    x    1     ?   0   0   1    0    ?  : ?  :  -;
      ?    *    ?     ?   0   0   1    0    ?  : 0  :  0;
      ?    x    ?     ?   0   0   1    0    ?  : 0  :  0;
      ?    x    ?     1   1   ?   1    0    ?  : 1  :  1;
      1    x    1     1   ?   ?   1    0    ?  : 1  :  1;
      ?    x    ?     0   1   ?   1    0    ?  : 0  :  0;
      ?    x    0     0   ?   ?   1    0    ?  : 0  :  1;
      0    x    ?     0   ?   ?   1    0    ?  : 0  :  0;
      ?    r    0     0   ?   ?   1    0    ?  : ?  :  1 ; 
      ?   (?0)  ?     ?   ?   ?   1    0    ?  : ?  :  -;  // no changes on falling clk edge
      1    r    1     ?   0   1   1    0    ?  : ?  :  1;
      0    r    ?     ?   0   1   1    0    ?  : ?  :  0;
      ?    r    0     ?   0   ?   1    0    ?  : ?  :  1;
      ?    x    0     ?   0   ?   1    0    ?  : 0  :  0;
      1    x    1     ?   0   ?   1    0    ?  : 1  :  1; // no changes when in switches
      0    x    ?     ?   0   ?   1    0    ?  : 0  :  0; // no changes when in switches
      1    *    1     ?   0   ?   1    0    ?  : 1  :  1; // reduce pessimism
      0    *    ?     ?   0   ?   1    0    ?  : 0  :  0; // reduce pessimism
      ?    ?    ?     ?   ?   ?   0    1    ?  : ?  :  x;
      ?    ?    ?     ?   ?   ?   1    1    ?  : ?  :  x;
      ?    ?    ?     ?   ?   ?   0    0    ?  : ?  :  x;

   endtable
endprimitive  // udp_sedffts 
*/

// $Id: udp_sedffsr.v
//
// verilog UDP for a 2-input mux used in scan cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//
 primitive udp_sedffsr_PWR (out, in, clk, clr_, set_, si, se, en, VDD, VSS, NOTIFIER);
   output out;  
   input  in, clk, clr_, set_, si, se,  en, VDD, VSS, NOTIFIER;
   reg    out;

   table
   // in  clk  clr_  set_ si  se  en  VDD   VSS   NOT : Qt : Qt+1
      ?    ?    ?     ?   ?   ?   ?   ?      ?     *  : ?  :  x; // any NOTIFIER changed
      ?    ?    0     1   ?   ?   ?   1      0     ?  : ?  :  0; 
      ?    ?    ?     0   ?   ?   ?   1      0     ?  : ?  :  1; 
      ?    r    ?     1   0   1   ?   1      0     ?  : ?  :  0;
      ?    r    1     ?   1   1   ?   1      0     ?  : ?  :  1;      
      ?    b    ?     1   ?   *   ?   1      0     ?  : 0  :  0; // no changes when se switches
      ?    b    1     ?   ?   *   ?   1      0     ?  : 1  :  1; // no changes when se switches
      ?    b    ?     1   *   ?   ?   1      0     ?  : 0  :  0; // no changes when si switches
      ?    b    1     ?   *   ?   ?   1      0     ?  : 1  :  1; // no changes when si switches
      *    b    ?     1   ?   ?   ?   1      0     ?  : 0  :  0; // no changes when in switches
      *    b    1     ?   ?   ?   ?   1      0     ?  : 1  :  1; // no changes when in switches
      ?    b    ?     1   ?   ?   *   1      0     ?  : 0  :  0; // no changes when en switches
      ?    b    1     ?   ?   ?   *   1      0     ?  : 1  :  1; // no changes when en switches
      ?    ?    *     1   ?   0   0   1      0     ?  : 0  :  0; //new
      ?    x    1     1   ?   0   0   1      0     ?  : 0  :  0;
      ?    x    1     1   ?   0   0   1      0     ?  : 1  :  1;
      ?    ?    *     1   0   ?   0   1      0     ?  : 0  :  0; //new
      0    ?    *     1   ?   0   1   1      0     ?  : 0  :  0; //new
      ?    b    *     1   ?   ?   ?   1      0     ?  : 0  :  0; //new
      ?    ?    1     *   ?   0   0   1      0     ?  : 1  :  1; //new
      ?    ?    1     *   1   ?   0   1      0     ?  : 1  :  1; //new
      1    ?    1     *   ?   0   1   1      0     ?  : 1  :  1; //new
      ?    b    1     *   ?   ?   ?   1      0     ?  : 1  :  1; //new
      ?    *    1     ?   1   1   ?   1      0     ?  : 1  :  1;
      ?    x    1     ?   1   1   ?   1      0     ?  : 1  :  1;
      ?    x    1     ?   ?   0   0   1      0     ?  : 1  :  1;
      ?    x    1     ?   1   ?   0   1      0     ?  : 1  :  1;
      ?    *    1     ?   1   ?   0   1      0     ?  : 1  :  1;
      ?    *    ?     1   0   1   ?   1      0     ?  : 0  :  0;
      ?    x    ?     1   0   1   ?   1      0     ?  : 0  :  0;
      ?    x    ?     1   ?   0   0   1      0     ?  : 0  :  0;
      ?    x    ?     1   0   ?   0   1      0     ?  : 0  :  0;
      ?    *    ?     1   0   ?   0   1      0     ?  : 0  :  0;
      0    r    ?     1   0   ?   1   1      0     ?  : ?  :  0 ; 
      0    *    ?     1   0   ?   ?   1      0     ?  : 0  :  0 ;
      0    x    ?     1   0   ?   ?   1      0     ?  : 0  :  0 ; 
      1    r    1     ?   1   ?   1   1      0     ?  : ?  :  1 ; 
      1    *    1     ?   1   ?   ?   1      0     ?  : 1  :  1 ; 
      1    x    1     ?   1   ?   ?   1      0     ?  : 1  :  1 ; 
      ?  (10)   ?     ?   ?   ?   ?   1      0     ?  : ?  :  -;  // no changes on falling clk edge
      ?  (x0)   ?     ?   ?   ?   ?   1      0     ?  : ?  :  -;  // no changes on falling clk edge
      1    r    1     ?   ?   0   1   1      0     ?  : ?  :  1;
      0    r    ?     1   ?   0   1   1      0     ?  : ?  :  0 ; 
      ?    *    ?     1   ?   0   0   1      0     ?  : 0  :  0;
      ?    *    1     ?   ?   0   0   1      0     ?  : 1  :  1;
      1    x    1     ?   ?   0   ?   1      0     ?  : 1  :  1; // no changes when in switches
      0    x    ?     1   ?   0   ?   1      0     ?  : 0  :  0; // no changes when in switches
      1    *    1     ?   ?   0   ?   1      0     ?  : 1  :  1; // reduce pessimism
      0    *    ?     1   ?   0   ?   1      0     ?  : 0  :  0; // reduce pessimism
      ?    ?    ?     ?   ?   ?   ?   0      1     ?  : ?  :  x; 
      ?    ?    ?     ?   ?   ?   ?   1      1     ?  : ?  :  x; 
      ?    ?    ?     ?   ?   ?   ?   0      0     ?  : ?  :  x; 

   endtable
endprimitive // udp_sedffsr
   
// $Id: udp_mux.v
//
// verilog UDP for a 2-input mux used in scan cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_mux_PWR (out, in, s_in, s_sel, VDD, VSS);
   output out;  
   input  in, s_in, s_sel, VDD, VSS;

   table

// in  s_in  s_sel VDD VSS :  out
//
   1  ?   0  1  0  :  1 ;
   0  ?   0  1  0  :  0 ;
   ?  1   1  1  0  :  1 ;
   ?  0   1  1  0  :  0 ;
   0  0   x  1  0  :  0 ;
   1  1   x  1  0  :  1 ;
   ?  ?   ?  0  1  :  x ;
   ?  ?   ?  1  1  :  x ;
   ?  ?   ?  0  0  :  x ;
   endtable
endprimitive // udp_mux

// $Id: udp_mux2.v
//
// verilog UDP for 2-input muxes
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_mux2_PWR (out, in0, in1, sel, VDD, VSS);
   output out;  
   input  in0, in1, sel, VDD, VSS;

   table

// in0 in1  sel VDD VSS :  out
//
   1  ?   0  1  0  :  1 ;
   0  ?   0  1  0  :  0 ;
   ?  1   1  1  0  :  1 ;
   ?  0   1  1  0  :  0 ;
   0  0   x  1  0  :  0 ;
   1  1   x  1  0  :  1 ;
   ?  ?   ?  0  0  :  x ;
   ?  ?   ?  0  1  :  x ;
   ?  ?   ?  1  1  :  x ;

   endtable
endprimitive // udp_mux2

// $Id: udp_mux4.v
//
// verilog UDP for 4-input muxes
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_mux4_PWR (out, in0, in1, in2, in3, sel_0, sel_1, VDD, VSS);
   output out;  
   input  in0, in1, in2, in3, sel_0, sel_1, VDD, VSS;

   table

// in0 in1 in2 in3 sel_0 sel_1 VDD VSS:  out
//
   0  ?  ?  ?  0  0  1  0  :  0;
   1  ?  ?  ?  0  0  1  0  :  1;
   ?  0  ?  ?  1  0  1  0  :  0;
   ?  1  ?  ?  1  0  1  0  :  1;
   ?  ?  0  ?  0  1  1  0  :  0;
   ?  ?  1  ?  0  1  1  0  :  1;
   ?  ?  ?  0  1  1  1  0  :  0;
   ?  ?  ?  1  1  1  1  0  :  1;
   0  0  ?  ?  x  0  1  0  :  0;
   1  1  ?  ?  x  0  1  0  :  1;
   ?  ?  0  0  x  1  1  0  :  0;
   ?  ?  1  1  x  1  1  0  :  1;
   0  ?  0  ?  0  x  1  0  :  0;
   1  ?  1  ?  0  x  1  0  :  1;
   ?  0  ?  0  1  x  1  0  :  0;
   ?  1  ?  1  1  x  1  0  :  1;
   1  1  1  1  x  x  1  0  :  1;
   0  0  0  0  x  x  1  0  :  0;
   ?  ?  ?  ?  ?  ?  0  0  :  x;
   ?  ?  ?  ?  ?  ?  0  1  :  x;
   ?  ?  ?  ?  ?  ?  1  1  :  x;

   endtable
endprimitive // udp_mux4

// $Id: udp_rslatn_out.v
//
// verilog UDP for the true output of rslatn cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_rslatn_out_PWR (out, r_, s_, VDD, VSS, NOTIFIER);
   output out;  
   input  r_, s_, VDD, VSS, NOTIFIER;
   reg    out;

   table

// r_  s_  VDD  VSS  NOT : Qt : Qt+1
// 
  (?1) 1   1   0   ?   : ?  :  -  ; // no change
   1  (?1) 1   0   ?   : ?  :  -  ; // no change
  (?0) 1   1   0   ?   : ?  :  0  ; // reset
   0  (?1) 1   0   ?   : ?  :  0  ; // reset
   ?   0   1   0   ?   : ?  :  1  ; // unused state
  (?1) x   1   0   ?   : 1  :  1  ; // reduced pessimism
   1  (?x) 1   0   ?   : 1  :  1  ; // reduced pessimism
  (?x) 1   1   0   ?   : 0  :  0  ; // reduced pessimism
   x  (?1) 1   0   ?   : 0  :  0  ; // reduced pessimism
   ?   ?   0   1   ?   : ?  :  x  ; 
   ?   ?   0   0   ?   : ?  :  x  ; 
   ?   ?   1   1   ?   : ?  :  x  ; 
   ?   ?   ?   ?   *   : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_rslatn_out

// $Id: udp_rslatn_out_.v
//
// verilog UDP for the complementary output of rslatn cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_rslatn_out__PWR (out_, r_, s_, VDD, VSS, NOTIFIER);
   output out_;  
   input  r_, s_, VDD, VSS, NOTIFIER;
   reg    out_;

   table

// r_  s_  VDD  VSS  NOT : Qt : Qt+1
// 
  (?1) 1   1   0    ?   : ?  :  -  ; // no change
   1  (?1) 1   0    ?   : ?  :  -  ; // no change
   0   ?   1   0    ?   : ?  :  1  ; // reset
  (?1) 0   1   0    ?   : ?  :  0  ; // set
   1  (?0) 1   0    ?   : ?  :  0  ; // set
  (?1) x   1   0    ?   : 0  :  0  ; // reduced pessimism
   1  (?x) 1   0    ?   : 0  :  0  ; // reduced pessimism
  (?x) 1   1   0    ?   : 1  :  1  ; // reduced pessimism
   x  (?1) 1   0    ?   : 1  :  1  ; // reduced pessimism
   ?   ?   0   0    ?   : ?  :  x  ; 
   ?   ?   0   1    ?   : ?  :  x  ; 
   ?   ?   1   1    ?   : ?  :  x  ; 
   ?   ?   ?   ?    *   : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_rslatn_out_

// $Id: udp_rslat_out.v
//
// verilog UDP for true output of rslat cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_rslat_out_PWR (out, r, s, VDD, VSS, NOTIFIER);
   output out;  
   input  r, s, VDD, VSS, NOTIFIER;
   reg    out;

   table

// r   s   VDD  VSS  NOT : Qt : Qt+1
// 
  (?0) 0   1   0   ?   : ?  :  -  ; // no change
   0  (?0) 1   0   ?   : ?  :  -  ; // no change
   1   ?   1   0   ?   : ?  :  0  ; // reset
  (?0) 1   1   0   ?   : ?  :  1  ; // set
   0  (?1) 1   0   ?   : ?  :  1  ; // set
  (?0) x   1   0   ?   : 1  :  1  ; // reduced pessimism
   0  (?x) 1   0   ?   : 1  :  1  ; // reduced pessimism
  (?x) 0   1   0   ?   : 0  :  0  ; // reduced pessimism
   x  (?0) 1   0   ?   : 0  :  0  ; // reduced pessimism
   ?   ?   0   1   ?   : ?  :  x  ;
   ?   ?   0   0   ?   : ?  :  x  ;
   ?   ?   1   1   ?   : ?  :  x  ;
   ?   ?   ?   ?   *   : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_rslat_out

// $Id: udp_rslat_out_.v
//
// verilog UDP for complementary output on rslat cells
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_rslat_out__PWR (out_, r, s, VDD, VSS, NOTIFIER);
   output out_;  
   input  r, s, VDD, VSS, NOTIFIER;
   reg    out_;

   table

// r   s   VDD  VSS  NOT : Qt : Qt+1
// 
  (?0) 0   1   0   ?   : ?  :  -  ; // no change
   0  (?0) 1   0   ?   : ?  :  -  ; // no change
  (?1) 0   1   0   ?   : ?  :  1  ; // reset
   1  (?0) 1   0   ?   : ?  :  1  ; // reset
   ?   1   1   0   ?   : ?  :  0  ; // set
  (?0) x   1   0   ?   : 0  :  0  ; // reduced pessimism
   0  (?x) 1   0   ?   : 0  :  0  ; // reduced pessimism
  (?x) 0   1   0   ?   : 1  :  1  ; // reduced pessimism
   x  (?0) 1   0   ?   : 1  :  1  ; // reduced pessimism
   ?   ?   0   0   ?   : ?  :  x  ; 
   ?   ?   0   1   ?   : ?  :  x  ; 
   ?   ?   1   1   ?   : ?  :  x  ; 
   ?   ?   ?   ?   *   : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_rslat_out_

// $Id: udp_tlat.v
//
// verilog UDP for d latches
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_tlat_PWR (out, in, hold, clr_, set_, VDD, VSS, NOTIFIER);
   output out;  
   input  in, hold, clr_, set_, VDD, VSS, NOTIFIER;
   reg    out;

   table

// in  hold  clr_   set_  VDD, VSS, NOT  : Qt : Qt+1
//
   1  0   1   ?   1   0   ?   : ?  :  1  ; // 
   0  0   ?   1   1   0   ?   : ?  :  0  ; // 
   1  *   1   ?   1   0   ?   : 1  :  1  ; // reduce pessimism
   0  *   ?   1   1   0   ?   : 0  :  0  ; // reduce pessimism
   *  1   ?   ?   1   0   ?   : ?  :  -  ; // no changes when in switches
   ?  ?   ?   0   1   0   ?   : ?  :  1  ; // set output
   ?  1   1   *   1   0   ?   : 1  :  1  ; // cover all transistions on set_
   1  ?   1   *   1   0   ?   : 1  :  1  ; // cover all transistions on set_
   ?  ?   0   1   1   0   ?   : ?  :  0  ; // reset output
   ?  1   *   1   1   0   ?   : 0  :  0  ; // cover all transistions on clr_
   0  ?   *   1   1   0   ?   : 0  :  0  ; // cover all transistions on clr_
   ?  ?   ?   ?   0   0   ?   : ?  :  x  ;
   ?  ?   ?   ?   0   1   ?   : ?  :  x  ;
   ?  ?   ?   ?   1   1   ?   : ?  :  x  ;
   ?  ?   ?   ?   ?   ?   *   : ?  :  x  ; // any NOTIFIER changed


   endtable
endprimitive // udp_tlat

//$Id udp_xgen.v
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_xgen_PWR (out, in, en, e, VDD, VSS);
   output out;  
   input  in, en, e, VDD, VSS;

   table

// in  en    e   VDD   VSS   : out;
//	     	  
   0   0     0    1    0     : x  ; // 
   0   0     1    1    0     : 0  ; // 
   0   1     0    1    0     : 0  ; // 
   0   1     1    1    0     : x  ; // 
   1   0     0    1    0     : x  ; // 
   1   0     1    1    0     : 1  ; // 
   1   1     0    1    0     : 1  ; // 
   1   1     1    1    0     : x  ; // 
   ?   ?     ?    0    0     : x  ; // 
   ?   ?     ?    0    1     : x  ; // 
   ?   ?     ?    1    1     : x  ; // 

   endtable
endprimitive // udp_xgen

//$Id udp_tlatrf.v
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_tlatrf_PWR (out, in, ww, wwn, VDD, VSS, NOTIFIER);
   output out;  
   input  in, ww, wwn, VDD, VSS, NOTIFIER;
   reg    out;

   table

// in  ww    wwn  VDD  VSS  NOT  : Qt : Qt+1
//	     
   1   ?     0    1	0	?    : ?  :  1  ; // 
   1   1     ?    1	0	?    : ?  :  1  ; // 
   0   ?     0    1	0	?    : ?  :  0  ; // 
   0   1     ?    1	0	?    : ?  :  0  ; // 
   1   *     ?    1	0	?    : 1  :  1  ; // reduce pessimism
   1   ?     *    1	0	?    : 1  :  1  ; // reduce pessimism
   0   *     ?    1	0	?    : 0  :  0  ; // reduce pessimism
   0   ?     *    1	0	?    : 0  :  0  ; // reduce pessimism
   *   0     1    1	0	?    : ?  :  -  ; // no changes when in switches
   ?   ?     ?    0	0	?    : ?  :  x  ; 
   ?   ?     ?    0	1	?    : ?  :  x  ; 
   ?   ?     ?    1	1	?    : ?  :  x  ; 
   ?   ?     ?    ?	?	*    : ?  :  x  ; // any NOTIFIER changed

   endtable
endprimitive // udp_tlatrf

//$Id udp_tlatrf2.v
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_tlatrf2_PWR (out, in1, w1w, in2, w2w, VDD, VSS, NOTIFIER);
   output out;  
   input  in1, w1w, VDD, VSS, NOTIFIER;
   input  in2, w2w;
   reg    out;

   table

// in1 ww1 in2 ww2  VDD  VSS  NOT  : Qt : Qt+1
//	     
   ?   ?    ?   ?    ?    ?   *    : ?  :  x  ; //
   1   1    ?   0    1    0   ?    : ?  :  1  ; //
   1   *    ?   0    1    0   ?    : 1  :  1  ; //
   0   1    ?   0    1    0   ?    : ?  :  0  ; //
   0   *    ?   0    1    0   ?    : 0  :  0  ; //
   ?   0    1   1    1    0   ?    : ?  :  1  ; //
   ?   0    1   *    1    0   ?    : 1  :  1  ; //
   ?   0    0   1    1    0   ?    : ?  :  0  ; //
   ?   0    0   *    1    0   ?    : 0  :  0  ; //
   *   0    ?   0    1    0   ?    : ?  :  -  ; //
   ?   0    *   0    1    0   ?    : ?  :  -  ; //
   1   *    1   1    1    0   ?    : ?  :  1  ; //
   1   1    1   *    1    0   ?    : ?  :  1  ; //
   0   *    0   1    1    0   ?    : ?  :  0  ; //
   0   1    0   *    1    0   ?    : ?  :  0  ; //
   ?   ?    ?   ?    0    0   ?    : ?  :  x  ;
   ?   ?    ?   ?    0    1   ?    : ?  :  x  ;
   ?   ?    ?   ?    1    1   ?    : ?  :  x  ;


   endtable
endprimitive // udp_tlatrf2

//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_outrf_PWR (out, in, rwn, rw, VDD, VSS);
   output out;  
   input  in, rwn, rw, VDD, VSS;

   table

// in  rwn   rw   VDD  VSS  : out;
//	     	  
   0   0     ?    1    0    : 1  ; // 
   1   ?     1    1    0    : 1  ; // 
   ?   1     0    1    0    : 0  ; // 
   1   ?     0    1    0    : 0  ; // 
   0   1     ?    1    0    : 0  ; // 
   ?   ?     ?    0    0    : x  ;
   ?   ?     ?    0    1    : x  ;
   ?   ?     ?    1    1    : x  ;

   endtable
endprimitive // udp_outrf

//$Id udp_bmx.v
//
// verilog UDP for 4-input muxes
//
//
// Library Service Department
// Design Service Division, SMIC
// Zhangjiang Rd.,Pudong New Area , Shanghai, PR of China 201203 
// (+8621)50802000
//
//
//

primitive udp_bmx_PWR (out, x2, a, s, m1, m0, VDD, VSS);
   output out;  
   input   x2, a, s, m1, m0, VDD, VSS;

   table

// x2 a  s m1 m0 VDD  VSS  :  out
//
   0  1  1  ?  ? 1    0    :  0;
   0  1  0  0  ? 1    0    :  1;
   0  1  0  1  ? 1    0    :  0;
   0  0  1  0  ? 1    0    :  0;
   0  0  1  1  ? 1    0    :  1;
   0  0  0  ?  ? 1    0    :  1;
   1  1  1  ?  ? 1    0    :  0;
   1  1  0  ?  0 1    0    :  1;
   1  1  0  ?  1 1    0    :  0;
   1  0  1  ?  0 1    0    :  0;
   1  0  1  ?  1 1    0    :  1;
   1  0  0  ?  ? 1    0    :  1;
   ?  ?  ?  ?  ? 0    0    :  x;
   ?  ?  ?  ?  ? 0    1    :  x;
   ?  ?  ?  ?  ? 1    1    :  x;

   endtable
endprimitive // udp_bmx
